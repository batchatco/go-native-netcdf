netcdf testvlen {
types:
  int(*) vint;

dimensions:
  dim = 6;

variables:
  vint v(dim);
  vint v2(dim);

data:
  v = {}, {1}, {2,3}, {4,5,6}, {7,8,9,10}, {11,12,13,14,15};
  v2 = {11,12,13,14,15}, {7,8,9,10}, {4,5,6}, {2,3}, {1}, {};
}
