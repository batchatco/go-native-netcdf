netcdf testtypes {
 dimensions:
  dim = 1;
  d1 = 2;
  d2 = 2;

 variables:
  int i32x2(d1, d2);

 data:
  i32x2 = -10000000, 10000000, -20000000, 20000000;
}
