netcdf testfills2 {
dimensions:
  dim = 1;
  d1 = 2;
  d2 = 2;
variables:
  string str;
  string str:_FillValue = "#";
  string strx1(dim);
  string strx1:_FillValue = "#";
  string strx2(d1, d2);
  string strx2:_FillValue = "#";
  float f32;
  f32:_FillValue = 0;
  float f32x1(dim);
  f32x1:_FillValue = 0;
  float f32x2(d1, d2);
  f32x2:_FillValue = 0;
  double f64;
  f64:_FillValue = 0;
  double f64x1(dim);
  f64x1:_FillValue = 0;
  double f64x2(d1, d2);
  f64x2:_FillValue = 0;
  byte i8;
  i8:_FillValue = 0;
  byte i8x1(dim);
  i8x1:_FillValue = 0;
  byte i8x2(d1, d2);
  i8x2:_FillValue = 0;
  ubyte ui8;
  ui8:_FillValue = 0;
  ubyte ui8x1(dim);
  ui8x1:_FillValue = 0;
  ubyte ui8x2(d1, d2);
  ui8x2:_FillValue = 0;
  short i16;
  i16:_FillValue = 0;
  short i16x1(dim);
  i16x1:_FillValue = 0;
  short i16x2(d1, d2);
  i16x2:_FillValue = 0;
  ushort ui16;
  ui16:_FillValue = 0;
  ushort ui16x1(dim);
  ui16x1:_FillValue = 0;
  ushort ui16x2(d1, d2);
  ui16x2:_FillValue = 0;
  int i32;
  i32:_FillValue = 0;
  int i32x1(dim);
  i32x1:_FillValue = 0;
  int i32x2(d1, d2);
  i32x2:_FillValue = 0;
  uint ui32;
  ui32:_FillValue = 0;
  uint ui32x1(dim);
  ui32x1:_FillValue = 0;
  uint ui32x2(d1, d2);
  ui32x2:_FillValue = 0;
  int64 i64;
  i64:_FillValue = 0;
  int64 i64x1(dim);
  i64x1:_FillValue = 0;
  int64 i64x2(d1, d2);
  i64x2:_FillValue = 0;
  uint64 ui64;
  ui64:_FillValue = 0;
  uint64 ui64x1(dim);
  ui64x1:_FillValue = 0;
  uint64 ui64x2(d1, d2);
  ui64x2:_FillValue = 0;
}
