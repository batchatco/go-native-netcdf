netcdf t2_modified {
dimensions:
	valid_time = 8760 ;
	pressure_level = 6 ;
	latitude = 37 ;
	longitude = 41 ;
variables:
	int64 number ;
		number:long_name = "ensemble member numerical id" ;
		number:units = "1" ;
		number:standard_name = "realization" ;
	int64 valid_time(valid_time) ;
		valid_time:long_name = "time" ;
		valid_time:standard_name = "time" ;
		valid_time:units = "seconds since 1970-01-01" ;
		valid_time:calendar = "proleptic_gregorian" ;
	double pressure_level(pressure_level) ;
		pressure_level:_FillValue = NaN ;
		pressure_level:long_name = "pressure" ;
		pressure_level:units = "hPa" ;
		pressure_level:positive = "down" ;
		pressure_level:stored_direction = "decreasing" ;
		pressure_level:standard_name = "air_pressure" ;
	double latitude(latitude) ;
		latitude:_FillValue = NaN ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:stored_direction = "decreasing" ;
	double longitude(longitude) ;
		longitude:_FillValue = NaN ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
	string expver(valid_time) ;

// global attributes:
		:GRIB_centre = "ecmf" ;
		:GRIB_centreDescription = "European Centre for Medium-Range Weather Forecasts" ;
		:GRIB_subCentre = 0LL ;
		:Conventions = "CF-1.7" ;
		:institution = "European Centre for Medium-Range Weather Forecasts" ;
		:history = "2024-11-18T12:20 GRIB to CDM+CF via cfgrib-0.9.14.1/ecCodes-2.36.0 with {\"source\": \"data.grib\", \"filter_by_keys\": {\"stream\": [\"oper\"]}, \"encode_cf\": [\"parameter\", \"time\", \"geography\", \"vertical\"]}" ;
data:

 number = 0 ;

 valid_time = 1640995200, 1640998800, 1641002400, 1641006000, 1641009600, 
    1641013200, 1641016800, 1641020400, 1641024000, 1641027600, 1641031200, 
    1641034800, 1641038400, 1641042000, 1641045600, 1641049200, 1641052800, 
    1641056400, 1641060000, 1641063600, 1641067200, 1641070800, 1641074400, 
    1641078000, 1641081600, 1641085200, 1641088800, 1641092400, 1641096000, 
    1641099600, 1641103200, 1641106800, 1641110400, 1641114000, 1641117600, 
    1641121200, 1641124800, 1641128400, 1641132000, 1641135600, 1641139200, 
    1641142800, 1641146400, 1641150000, 1641153600, 1641157200, 1641160800, 
    1641164400, 1641168000, 1641171600, 1641175200, 1641178800, 1641182400, 
    1641186000, 1641189600, 1641193200, 1641196800, 1641200400, 1641204000, 
    1641207600, 1641211200, 1641214800, 1641218400, 1641222000, 1641225600, 
    1641229200, 1641232800, 1641236400, 1641240000, 1641243600, 1641247200, 
    1641250800, 1641254400, 1641258000, 1641261600, 1641265200, 1641268800, 
    1641272400, 1641276000, 1641279600, 1641283200, 1641286800, 1641290400, 
    1641294000, 1641297600, 1641301200, 1641304800, 1641308400, 1641312000, 
    1641315600, 1641319200, 1641322800, 1641326400, 1641330000, 1641333600, 
    1641337200, 1641340800, 1641344400, 1641348000, 1641351600, 1641355200, 
    1641358800, 1641362400, 1641366000, 1641369600, 1641373200, 1641376800, 
    1641380400, 1641384000, 1641387600, 1641391200, 1641394800, 1641398400, 
    1641402000, 1641405600, 1641409200, 1641412800, 1641416400, 1641420000, 
    1641423600, 1641427200, 1641430800, 1641434400, 1641438000, 1641441600, 
    1641445200, 1641448800, 1641452400, 1641456000, 1641459600, 1641463200, 
    1641466800, 1641470400, 1641474000, 1641477600, 1641481200, 1641484800, 
    1641488400, 1641492000, 1641495600, 1641499200, 1641502800, 1641506400, 
    1641510000, 1641513600, 1641517200, 1641520800, 1641524400, 1641528000, 
    1641531600, 1641535200, 1641538800, 1641542400, 1641546000, 1641549600, 
    1641553200, 1641556800, 1641560400, 1641564000, 1641567600, 1641571200, 
    1641574800, 1641578400, 1641582000, 1641585600, 1641589200, 1641592800, 
    1641596400, 1641600000, 1641603600, 1641607200, 1641610800, 1641614400, 
    1641618000, 1641621600, 1641625200, 1641628800, 1641632400, 1641636000, 
    1641639600, 1641643200, 1641646800, 1641650400, 1641654000, 1641657600, 
    1641661200, 1641664800, 1641668400, 1641672000, 1641675600, 1641679200, 
    1641682800, 1641686400, 1641690000, 1641693600, 1641697200, 1641700800, 
    1641704400, 1641708000, 1641711600, 1641715200, 1641718800, 1641722400, 
    1641726000, 1641729600, 1641733200, 1641736800, 1641740400, 1641744000, 
    1641747600, 1641751200, 1641754800, 1641758400, 1641762000, 1641765600, 
    1641769200, 1641772800, 1641776400, 1641780000, 1641783600, 1641787200, 
    1641790800, 1641794400, 1641798000, 1641801600, 1641805200, 1641808800, 
    1641812400, 1641816000, 1641819600, 1641823200, 1641826800, 1641830400, 
    1641834000, 1641837600, 1641841200, 1641844800, 1641848400, 1641852000, 
    1641855600, 1641859200, 1641862800, 1641866400, 1641870000, 1641873600, 
    1641877200, 1641880800, 1641884400, 1641888000, 1641891600, 1641895200, 
    1641898800, 1641902400, 1641906000, 1641909600, 1641913200, 1641916800, 
    1641920400, 1641924000, 1641927600, 1641931200, 1641934800, 1641938400, 
    1641942000, 1641945600, 1641949200, 1641952800, 1641956400, 1641960000, 
    1641963600, 1641967200, 1641970800, 1641974400, 1641978000, 1641981600, 
    1641985200, 1641988800, 1641992400, 1641996000, 1641999600, 1642003200, 
    1642006800, 1642010400, 1642014000, 1642017600, 1642021200, 1642024800, 
    1642028400, 1642032000, 1642035600, 1642039200, 1642042800, 1642046400, 
    1642050000, 1642053600, 1642057200, 1642060800, 1642064400, 1642068000, 
    1642071600, 1642075200, 1642078800, 1642082400, 1642086000, 1642089600, 
    1642093200, 1642096800, 1642100400, 1642104000, 1642107600, 1642111200, 
    1642114800, 1642118400, 1642122000, 1642125600, 1642129200, 1642132800, 
    1642136400, 1642140000, 1642143600, 1642147200, 1642150800, 1642154400, 
    1642158000, 1642161600, 1642165200, 1642168800, 1642172400, 1642176000, 
    1642179600, 1642183200, 1642186800, 1642190400, 1642194000, 1642197600, 
    1642201200, 1642204800, 1642208400, 1642212000, 1642215600, 1642219200, 
    1642222800, 1642226400, 1642230000, 1642233600, 1642237200, 1642240800, 
    1642244400, 1642248000, 1642251600, 1642255200, 1642258800, 1642262400, 
    1642266000, 1642269600, 1642273200, 1642276800, 1642280400, 1642284000, 
    1642287600, 1642291200, 1642294800, 1642298400, 1642302000, 1642305600, 
    1642309200, 1642312800, 1642316400, 1642320000, 1642323600, 1642327200, 
    1642330800, 1642334400, 1642338000, 1642341600, 1642345200, 1642348800, 
    1642352400, 1642356000, 1642359600, 1642363200, 1642366800, 1642370400, 
    1642374000, 1642377600, 1642381200, 1642384800, 1642388400, 1642392000, 
    1642395600, 1642399200, 1642402800, 1642406400, 1642410000, 1642413600, 
    1642417200, 1642420800, 1642424400, 1642428000, 1642431600, 1642435200, 
    1642438800, 1642442400, 1642446000, 1642449600, 1642453200, 1642456800, 
    1642460400, 1642464000, 1642467600, 1642471200, 1642474800, 1642478400, 
    1642482000, 1642485600, 1642489200, 1642492800, 1642496400, 1642500000, 
    1642503600, 1642507200, 1642510800, 1642514400, 1642518000, 1642521600, 
    1642525200, 1642528800, 1642532400, 1642536000, 1642539600, 1642543200, 
    1642546800, 1642550400, 1642554000, 1642557600, 1642561200, 1642564800, 
    1642568400, 1642572000, 1642575600, 1642579200, 1642582800, 1642586400, 
    1642590000, 1642593600, 1642597200, 1642600800, 1642604400, 1642608000, 
    1642611600, 1642615200, 1642618800, 1642622400, 1642626000, 1642629600, 
    1642633200, 1642636800, 1642640400, 1642644000, 1642647600, 1642651200, 
    1642654800, 1642658400, 1642662000, 1642665600, 1642669200, 1642672800, 
    1642676400, 1642680000, 1642683600, 1642687200, 1642690800, 1642694400, 
    1642698000, 1642701600, 1642705200, 1642708800, 1642712400, 1642716000, 
    1642719600, 1642723200, 1642726800, 1642730400, 1642734000, 1642737600, 
    1642741200, 1642744800, 1642748400, 1642752000, 1642755600, 1642759200, 
    1642762800, 1642766400, 1642770000, 1642773600, 1642777200, 1642780800, 
    1642784400, 1642788000, 1642791600, 1642795200, 1642798800, 1642802400, 
    1642806000, 1642809600, 1642813200, 1642816800, 1642820400, 1642824000, 
    1642827600, 1642831200, 1642834800, 1642838400, 1642842000, 1642845600, 
    1642849200, 1642852800, 1642856400, 1642860000, 1642863600, 1642867200, 
    1642870800, 1642874400, 1642878000, 1642881600, 1642885200, 1642888800, 
    1642892400, 1642896000, 1642899600, 1642903200, 1642906800, 1642910400, 
    1642914000, 1642917600, 1642921200, 1642924800, 1642928400, 1642932000, 
    1642935600, 1642939200, 1642942800, 1642946400, 1642950000, 1642953600, 
    1642957200, 1642960800, 1642964400, 1642968000, 1642971600, 1642975200, 
    1642978800, 1642982400, 1642986000, 1642989600, 1642993200, 1642996800, 
    1643000400, 1643004000, 1643007600, 1643011200, 1643014800, 1643018400, 
    1643022000, 1643025600, 1643029200, 1643032800, 1643036400, 1643040000, 
    1643043600, 1643047200, 1643050800, 1643054400, 1643058000, 1643061600, 
    1643065200, 1643068800, 1643072400, 1643076000, 1643079600, 1643083200, 
    1643086800, 1643090400, 1643094000, 1643097600, 1643101200, 1643104800, 
    1643108400, 1643112000, 1643115600, 1643119200, 1643122800, 1643126400, 
    1643130000, 1643133600, 1643137200, 1643140800, 1643144400, 1643148000, 
    1643151600, 1643155200, 1643158800, 1643162400, 1643166000, 1643169600, 
    1643173200, 1643176800, 1643180400, 1643184000, 1643187600, 1643191200, 
    1643194800, 1643198400, 1643202000, 1643205600, 1643209200, 1643212800, 
    1643216400, 1643220000, 1643223600, 1643227200, 1643230800, 1643234400, 
    1643238000, 1643241600, 1643245200, 1643248800, 1643252400, 1643256000, 
    1643259600, 1643263200, 1643266800, 1643270400, 1643274000, 1643277600, 
    1643281200, 1643284800, 1643288400, 1643292000, 1643295600, 1643299200, 
    1643302800, 1643306400, 1643310000, 1643313600, 1643317200, 1643320800, 
    1643324400, 1643328000, 1643331600, 1643335200, 1643338800, 1643342400, 
    1643346000, 1643349600, 1643353200, 1643356800, 1643360400, 1643364000, 
    1643367600, 1643371200, 1643374800, 1643378400, 1643382000, 1643385600, 
    1643389200, 1643392800, 1643396400, 1643400000, 1643403600, 1643407200, 
    1643410800, 1643414400, 1643418000, 1643421600, 1643425200, 1643428800, 
    1643432400, 1643436000, 1643439600, 1643443200, 1643446800, 1643450400, 
    1643454000, 1643457600, 1643461200, 1643464800, 1643468400, 1643472000, 
    1643475600, 1643479200, 1643482800, 1643486400, 1643490000, 1643493600, 
    1643497200, 1643500800, 1643504400, 1643508000, 1643511600, 1643515200, 
    1643518800, 1643522400, 1643526000, 1643529600, 1643533200, 1643536800, 
    1643540400, 1643544000, 1643547600, 1643551200, 1643554800, 1643558400, 
    1643562000, 1643565600, 1643569200, 1643572800, 1643576400, 1643580000, 
    1643583600, 1643587200, 1643590800, 1643594400, 1643598000, 1643601600, 
    1643605200, 1643608800, 1643612400, 1643616000, 1643619600, 1643623200, 
    1643626800, 1643630400, 1643634000, 1643637600, 1643641200, 1643644800, 
    1643648400, 1643652000, 1643655600, 1643659200, 1643662800, 1643666400, 
    1643670000, 1643673600, 1643677200, 1643680800, 1643684400, 1643688000, 
    1643691600, 1643695200, 1643698800, 1643702400, 1643706000, 1643709600, 
    1643713200, 1643716800, 1643720400, 1643724000, 1643727600, 1643731200, 
    1643734800, 1643738400, 1643742000, 1643745600, 1643749200, 1643752800, 
    1643756400, 1643760000, 1643763600, 1643767200, 1643770800, 1643774400, 
    1643778000, 1643781600, 1643785200, 1643788800, 1643792400, 1643796000, 
    1643799600, 1643803200, 1643806800, 1643810400, 1643814000, 1643817600, 
    1643821200, 1643824800, 1643828400, 1643832000, 1643835600, 1643839200, 
    1643842800, 1643846400, 1643850000, 1643853600, 1643857200, 1643860800, 
    1643864400, 1643868000, 1643871600, 1643875200, 1643878800, 1643882400, 
    1643886000, 1643889600, 1643893200, 1643896800, 1643900400, 1643904000, 
    1643907600, 1643911200, 1643914800, 1643918400, 1643922000, 1643925600, 
    1643929200, 1643932800, 1643936400, 1643940000, 1643943600, 1643947200, 
    1643950800, 1643954400, 1643958000, 1643961600, 1643965200, 1643968800, 
    1643972400, 1643976000, 1643979600, 1643983200, 1643986800, 1643990400, 
    1643994000, 1643997600, 1644001200, 1644004800, 1644008400, 1644012000, 
    1644015600, 1644019200, 1644022800, 1644026400, 1644030000, 1644033600, 
    1644037200, 1644040800, 1644044400, 1644048000, 1644051600, 1644055200, 
    1644058800, 1644062400, 1644066000, 1644069600, 1644073200, 1644076800, 
    1644080400, 1644084000, 1644087600, 1644091200, 1644094800, 1644098400, 
    1644102000, 1644105600, 1644109200, 1644112800, 1644116400, 1644120000, 
    1644123600, 1644127200, 1644130800, 1644134400, 1644138000, 1644141600, 
    1644145200, 1644148800, 1644152400, 1644156000, 1644159600, 1644163200, 
    1644166800, 1644170400, 1644174000, 1644177600, 1644181200, 1644184800, 
    1644188400, 1644192000, 1644195600, 1644199200, 1644202800, 1644206400, 
    1644210000, 1644213600, 1644217200, 1644220800, 1644224400, 1644228000, 
    1644231600, 1644235200, 1644238800, 1644242400, 1644246000, 1644249600, 
    1644253200, 1644256800, 1644260400, 1644264000, 1644267600, 1644271200, 
    1644274800, 1644278400, 1644282000, 1644285600, 1644289200, 1644292800, 
    1644296400, 1644300000, 1644303600, 1644307200, 1644310800, 1644314400, 
    1644318000, 1644321600, 1644325200, 1644328800, 1644332400, 1644336000, 
    1644339600, 1644343200, 1644346800, 1644350400, 1644354000, 1644357600, 
    1644361200, 1644364800, 1644368400, 1644372000, 1644375600, 1644379200, 
    1644382800, 1644386400, 1644390000, 1644393600, 1644397200, 1644400800, 
    1644404400, 1644408000, 1644411600, 1644415200, 1644418800, 1644422400, 
    1644426000, 1644429600, 1644433200, 1644436800, 1644440400, 1644444000, 
    1644447600, 1644451200, 1644454800, 1644458400, 1644462000, 1644465600, 
    1644469200, 1644472800, 1644476400, 1644480000, 1644483600, 1644487200, 
    1644490800, 1644494400, 1644498000, 1644501600, 1644505200, 1644508800, 
    1644512400, 1644516000, 1644519600, 1644523200, 1644526800, 1644530400, 
    1644534000, 1644537600, 1644541200, 1644544800, 1644548400, 1644552000, 
    1644555600, 1644559200, 1644562800, 1644566400, 1644570000, 1644573600, 
    1644577200, 1644580800, 1644584400, 1644588000, 1644591600, 1644595200, 
    1644598800, 1644602400, 1644606000, 1644609600, 1644613200, 1644616800, 
    1644620400, 1644624000, 1644627600, 1644631200, 1644634800, 1644638400, 
    1644642000, 1644645600, 1644649200, 1644652800, 1644656400, 1644660000, 
    1644663600, 1644667200, 1644670800, 1644674400, 1644678000, 1644681600, 
    1644685200, 1644688800, 1644692400, 1644696000, 1644699600, 1644703200, 
    1644706800, 1644710400, 1644714000, 1644717600, 1644721200, 1644724800, 
    1644728400, 1644732000, 1644735600, 1644739200, 1644742800, 1644746400, 
    1644750000, 1644753600, 1644757200, 1644760800, 1644764400, 1644768000, 
    1644771600, 1644775200, 1644778800, 1644782400, 1644786000, 1644789600, 
    1644793200, 1644796800, 1644800400, 1644804000, 1644807600, 1644811200, 
    1644814800, 1644818400, 1644822000, 1644825600, 1644829200, 1644832800, 
    1644836400, 1644840000, 1644843600, 1644847200, 1644850800, 1644854400, 
    1644858000, 1644861600, 1644865200, 1644868800, 1644872400, 1644876000, 
    1644879600, 1644883200, 1644886800, 1644890400, 1644894000, 1644897600, 
    1644901200, 1644904800, 1644908400, 1644912000, 1644915600, 1644919200, 
    1644922800, 1644926400, 1644930000, 1644933600, 1644937200, 1644940800, 
    1644944400, 1644948000, 1644951600, 1644955200, 1644958800, 1644962400, 
    1644966000, 1644969600, 1644973200, 1644976800, 1644980400, 1644984000, 
    1644987600, 1644991200, 1644994800, 1644998400, 1645002000, 1645005600, 
    1645009200, 1645012800, 1645016400, 1645020000, 1645023600, 1645027200, 
    1645030800, 1645034400, 1645038000, 1645041600, 1645045200, 1645048800, 
    1645052400, 1645056000, 1645059600, 1645063200, 1645066800, 1645070400, 
    1645074000, 1645077600, 1645081200, 1645084800, 1645088400, 1645092000, 
    1645095600, 1645099200, 1645102800, 1645106400, 1645110000, 1645113600, 
    1645117200, 1645120800, 1645124400, 1645128000, 1645131600, 1645135200, 
    1645138800, 1645142400, 1645146000, 1645149600, 1645153200, 1645156800, 
    1645160400, 1645164000, 1645167600, 1645171200, 1645174800, 1645178400, 
    1645182000, 1645185600, 1645189200, 1645192800, 1645196400, 1645200000, 
    1645203600, 1645207200, 1645210800, 1645214400, 1645218000, 1645221600, 
    1645225200, 1645228800, 1645232400, 1645236000, 1645239600, 1645243200, 
    1645246800, 1645250400, 1645254000, 1645257600, 1645261200, 1645264800, 
    1645268400, 1645272000, 1645275600, 1645279200, 1645282800, 1645286400, 
    1645290000, 1645293600, 1645297200, 1645300800, 1645304400, 1645308000, 
    1645311600, 1645315200, 1645318800, 1645322400, 1645326000, 1645329600, 
    1645333200, 1645336800, 1645340400, 1645344000, 1645347600, 1645351200, 
    1645354800, 1645358400, 1645362000, 1645365600, 1645369200, 1645372800, 
    1645376400, 1645380000, 1645383600, 1645387200, 1645390800, 1645394400, 
    1645398000, 1645401600, 1645405200, 1645408800, 1645412400, 1645416000, 
    1645419600, 1645423200, 1645426800, 1645430400, 1645434000, 1645437600, 
    1645441200, 1645444800, 1645448400, 1645452000, 1645455600, 1645459200, 
    1645462800, 1645466400, 1645470000, 1645473600, 1645477200, 1645480800, 
    1645484400, 1645488000, 1645491600, 1645495200, 1645498800, 1645502400, 
    1645506000, 1645509600, 1645513200, 1645516800, 1645520400, 1645524000, 
    1645527600, 1645531200, 1645534800, 1645538400, 1645542000, 1645545600, 
    1645549200, 1645552800, 1645556400, 1645560000, 1645563600, 1645567200, 
    1645570800, 1645574400, 1645578000, 1645581600, 1645585200, 1645588800, 
    1645592400, 1645596000, 1645599600, 1645603200, 1645606800, 1645610400, 
    1645614000, 1645617600, 1645621200, 1645624800, 1645628400, 1645632000, 
    1645635600, 1645639200, 1645642800, 1645646400, 1645650000, 1645653600, 
    1645657200, 1645660800, 1645664400, 1645668000, 1645671600, 1645675200, 
    1645678800, 1645682400, 1645686000, 1645689600, 1645693200, 1645696800, 
    1645700400, 1645704000, 1645707600, 1645711200, 1645714800, 1645718400, 
    1645722000, 1645725600, 1645729200, 1645732800, 1645736400, 1645740000, 
    1645743600, 1645747200, 1645750800, 1645754400, 1645758000, 1645761600, 
    1645765200, 1645768800, 1645772400, 1645776000, 1645779600, 1645783200, 
    1645786800, 1645790400, 1645794000, 1645797600, 1645801200, 1645804800, 
    1645808400, 1645812000, 1645815600, 1645819200, 1645822800, 1645826400, 
    1645830000, 1645833600, 1645837200, 1645840800, 1645844400, 1645848000, 
    1645851600, 1645855200, 1645858800, 1645862400, 1645866000, 1645869600, 
    1645873200, 1645876800, 1645880400, 1645884000, 1645887600, 1645891200, 
    1645894800, 1645898400, 1645902000, 1645905600, 1645909200, 1645912800, 
    1645916400, 1645920000, 1645923600, 1645927200, 1645930800, 1645934400, 
    1645938000, 1645941600, 1645945200, 1645948800, 1645952400, 1645956000, 
    1645959600, 1645963200, 1645966800, 1645970400, 1645974000, 1645977600, 
    1645981200, 1645984800, 1645988400, 1645992000, 1645995600, 1645999200, 
    1646002800, 1646006400, 1646010000, 1646013600, 1646017200, 1646020800, 
    1646024400, 1646028000, 1646031600, 1646035200, 1646038800, 1646042400, 
    1646046000, 1646049600, 1646053200, 1646056800, 1646060400, 1646064000, 
    1646067600, 1646071200, 1646074800, 1646078400, 1646082000, 1646085600, 
    1646089200, 1646092800, 1646096400, 1646100000, 1646103600, 1646107200, 
    1646110800, 1646114400, 1646118000, 1646121600, 1646125200, 1646128800, 
    1646132400, 1646136000, 1646139600, 1646143200, 1646146800, 1646150400, 
    1646154000, 1646157600, 1646161200, 1646164800, 1646168400, 1646172000, 
    1646175600, 1646179200, 1646182800, 1646186400, 1646190000, 1646193600, 
    1646197200, 1646200800, 1646204400, 1646208000, 1646211600, 1646215200, 
    1646218800, 1646222400, 1646226000, 1646229600, 1646233200, 1646236800, 
    1646240400, 1646244000, 1646247600, 1646251200, 1646254800, 1646258400, 
    1646262000, 1646265600, 1646269200, 1646272800, 1646276400, 1646280000, 
    1646283600, 1646287200, 1646290800, 1646294400, 1646298000, 1646301600, 
    1646305200, 1646308800, 1646312400, 1646316000, 1646319600, 1646323200, 
    1646326800, 1646330400, 1646334000, 1646337600, 1646341200, 1646344800, 
    1646348400, 1646352000, 1646355600, 1646359200, 1646362800, 1646366400, 
    1646370000, 1646373600, 1646377200, 1646380800, 1646384400, 1646388000, 
    1646391600, 1646395200, 1646398800, 1646402400, 1646406000, 1646409600, 
    1646413200, 1646416800, 1646420400, 1646424000, 1646427600, 1646431200, 
    1646434800, 1646438400, 1646442000, 1646445600, 1646449200, 1646452800, 
    1646456400, 1646460000, 1646463600, 1646467200, 1646470800, 1646474400, 
    1646478000, 1646481600, 1646485200, 1646488800, 1646492400, 1646496000, 
    1646499600, 1646503200, 1646506800, 1646510400, 1646514000, 1646517600, 
    1646521200, 1646524800, 1646528400, 1646532000, 1646535600, 1646539200, 
    1646542800, 1646546400, 1646550000, 1646553600, 1646557200, 1646560800, 
    1646564400, 1646568000, 1646571600, 1646575200, 1646578800, 1646582400, 
    1646586000, 1646589600, 1646593200, 1646596800, 1646600400, 1646604000, 
    1646607600, 1646611200, 1646614800, 1646618400, 1646622000, 1646625600, 
    1646629200, 1646632800, 1646636400, 1646640000, 1646643600, 1646647200, 
    1646650800, 1646654400, 1646658000, 1646661600, 1646665200, 1646668800, 
    1646672400, 1646676000, 1646679600, 1646683200, 1646686800, 1646690400, 
    1646694000, 1646697600, 1646701200, 1646704800, 1646708400, 1646712000, 
    1646715600, 1646719200, 1646722800, 1646726400, 1646730000, 1646733600, 
    1646737200, 1646740800, 1646744400, 1646748000, 1646751600, 1646755200, 
    1646758800, 1646762400, 1646766000, 1646769600, 1646773200, 1646776800, 
    1646780400, 1646784000, 1646787600, 1646791200, 1646794800, 1646798400, 
    1646802000, 1646805600, 1646809200, 1646812800, 1646816400, 1646820000, 
    1646823600, 1646827200, 1646830800, 1646834400, 1646838000, 1646841600, 
    1646845200, 1646848800, 1646852400, 1646856000, 1646859600, 1646863200, 
    1646866800, 1646870400, 1646874000, 1646877600, 1646881200, 1646884800, 
    1646888400, 1646892000, 1646895600, 1646899200, 1646902800, 1646906400, 
    1646910000, 1646913600, 1646917200, 1646920800, 1646924400, 1646928000, 
    1646931600, 1646935200, 1646938800, 1646942400, 1646946000, 1646949600, 
    1646953200, 1646956800, 1646960400, 1646964000, 1646967600, 1646971200, 
    1646974800, 1646978400, 1646982000, 1646985600, 1646989200, 1646992800, 
    1646996400, 1647000000, 1647003600, 1647007200, 1647010800, 1647014400, 
    1647018000, 1647021600, 1647025200, 1647028800, 1647032400, 1647036000, 
    1647039600, 1647043200, 1647046800, 1647050400, 1647054000, 1647057600, 
    1647061200, 1647064800, 1647068400, 1647072000, 1647075600, 1647079200, 
    1647082800, 1647086400, 1647090000, 1647093600, 1647097200, 1647100800, 
    1647104400, 1647108000, 1647111600, 1647115200, 1647118800, 1647122400, 
    1647126000, 1647129600, 1647133200, 1647136800, 1647140400, 1647144000, 
    1647147600, 1647151200, 1647154800, 1647158400, 1647162000, 1647165600, 
    1647169200, 1647172800, 1647176400, 1647180000, 1647183600, 1647187200, 
    1647190800, 1647194400, 1647198000, 1647201600, 1647205200, 1647208800, 
    1647212400, 1647216000, 1647219600, 1647223200, 1647226800, 1647230400, 
    1647234000, 1647237600, 1647241200, 1647244800, 1647248400, 1647252000, 
    1647255600, 1647259200, 1647262800, 1647266400, 1647270000, 1647273600, 
    1647277200, 1647280800, 1647284400, 1647288000, 1647291600, 1647295200, 
    1647298800, 1647302400, 1647306000, 1647309600, 1647313200, 1647316800, 
    1647320400, 1647324000, 1647327600, 1647331200, 1647334800, 1647338400, 
    1647342000, 1647345600, 1647349200, 1647352800, 1647356400, 1647360000, 
    1647363600, 1647367200, 1647370800, 1647374400, 1647378000, 1647381600, 
    1647385200, 1647388800, 1647392400, 1647396000, 1647399600, 1647403200, 
    1647406800, 1647410400, 1647414000, 1647417600, 1647421200, 1647424800, 
    1647428400, 1647432000, 1647435600, 1647439200, 1647442800, 1647446400, 
    1647450000, 1647453600, 1647457200, 1647460800, 1647464400, 1647468000, 
    1647471600, 1647475200, 1647478800, 1647482400, 1647486000, 1647489600, 
    1647493200, 1647496800, 1647500400, 1647504000, 1647507600, 1647511200, 
    1647514800, 1647518400, 1647522000, 1647525600, 1647529200, 1647532800, 
    1647536400, 1647540000, 1647543600, 1647547200, 1647550800, 1647554400, 
    1647558000, 1647561600, 1647565200, 1647568800, 1647572400, 1647576000, 
    1647579600, 1647583200, 1647586800, 1647590400, 1647594000, 1647597600, 
    1647601200, 1647604800, 1647608400, 1647612000, 1647615600, 1647619200, 
    1647622800, 1647626400, 1647630000, 1647633600, 1647637200, 1647640800, 
    1647644400, 1647648000, 1647651600, 1647655200, 1647658800, 1647662400, 
    1647666000, 1647669600, 1647673200, 1647676800, 1647680400, 1647684000, 
    1647687600, 1647691200, 1647694800, 1647698400, 1647702000, 1647705600, 
    1647709200, 1647712800, 1647716400, 1647720000, 1647723600, 1647727200, 
    1647730800, 1647734400, 1647738000, 1647741600, 1647745200, 1647748800, 
    1647752400, 1647756000, 1647759600, 1647763200, 1647766800, 1647770400, 
    1647774000, 1647777600, 1647781200, 1647784800, 1647788400, 1647792000, 
    1647795600, 1647799200, 1647802800, 1647806400, 1647810000, 1647813600, 
    1647817200, 1647820800, 1647824400, 1647828000, 1647831600, 1647835200, 
    1647838800, 1647842400, 1647846000, 1647849600, 1647853200, 1647856800, 
    1647860400, 1647864000, 1647867600, 1647871200, 1647874800, 1647878400, 
    1647882000, 1647885600, 1647889200, 1647892800, 1647896400, 1647900000, 
    1647903600, 1647907200, 1647910800, 1647914400, 1647918000, 1647921600, 
    1647925200, 1647928800, 1647932400, 1647936000, 1647939600, 1647943200, 
    1647946800, 1647950400, 1647954000, 1647957600, 1647961200, 1647964800, 
    1647968400, 1647972000, 1647975600, 1647979200, 1647982800, 1647986400, 
    1647990000, 1647993600, 1647997200, 1648000800, 1648004400, 1648008000, 
    1648011600, 1648015200, 1648018800, 1648022400, 1648026000, 1648029600, 
    1648033200, 1648036800, 1648040400, 1648044000, 1648047600, 1648051200, 
    1648054800, 1648058400, 1648062000, 1648065600, 1648069200, 1648072800, 
    1648076400, 1648080000, 1648083600, 1648087200, 1648090800, 1648094400, 
    1648098000, 1648101600, 1648105200, 1648108800, 1648112400, 1648116000, 
    1648119600, 1648123200, 1648126800, 1648130400, 1648134000, 1648137600, 
    1648141200, 1648144800, 1648148400, 1648152000, 1648155600, 1648159200, 
    1648162800, 1648166400, 1648170000, 1648173600, 1648177200, 1648180800, 
    1648184400, 1648188000, 1648191600, 1648195200, 1648198800, 1648202400, 
    1648206000, 1648209600, 1648213200, 1648216800, 1648220400, 1648224000, 
    1648227600, 1648231200, 1648234800, 1648238400, 1648242000, 1648245600, 
    1648249200, 1648252800, 1648256400, 1648260000, 1648263600, 1648267200, 
    1648270800, 1648274400, 1648278000, 1648281600, 1648285200, 1648288800, 
    1648292400, 1648296000, 1648299600, 1648303200, 1648306800, 1648310400, 
    1648314000, 1648317600, 1648321200, 1648324800, 1648328400, 1648332000, 
    1648335600, 1648339200, 1648342800, 1648346400, 1648350000, 1648353600, 
    1648357200, 1648360800, 1648364400, 1648368000, 1648371600, 1648375200, 
    1648378800, 1648382400, 1648386000, 1648389600, 1648393200, 1648396800, 
    1648400400, 1648404000, 1648407600, 1648411200, 1648414800, 1648418400, 
    1648422000, 1648425600, 1648429200, 1648432800, 1648436400, 1648440000, 
    1648443600, 1648447200, 1648450800, 1648454400, 1648458000, 1648461600, 
    1648465200, 1648468800, 1648472400, 1648476000, 1648479600, 1648483200, 
    1648486800, 1648490400, 1648494000, 1648497600, 1648501200, 1648504800, 
    1648508400, 1648512000, 1648515600, 1648519200, 1648522800, 1648526400, 
    1648530000, 1648533600, 1648537200, 1648540800, 1648544400, 1648548000, 
    1648551600, 1648555200, 1648558800, 1648562400, 1648566000, 1648569600, 
    1648573200, 1648576800, 1648580400, 1648584000, 1648587600, 1648591200, 
    1648594800, 1648598400, 1648602000, 1648605600, 1648609200, 1648612800, 
    1648616400, 1648620000, 1648623600, 1648627200, 1648630800, 1648634400, 
    1648638000, 1648641600, 1648645200, 1648648800, 1648652400, 1648656000, 
    1648659600, 1648663200, 1648666800, 1648670400, 1648674000, 1648677600, 
    1648681200, 1648684800, 1648688400, 1648692000, 1648695600, 1648699200, 
    1648702800, 1648706400, 1648710000, 1648713600, 1648717200, 1648720800, 
    1648724400, 1648728000, 1648731600, 1648735200, 1648738800, 1648742400, 
    1648746000, 1648749600, 1648753200, 1648756800, 1648760400, 1648764000, 
    1648767600, 1648771200, 1648774800, 1648778400, 1648782000, 1648785600, 
    1648789200, 1648792800, 1648796400, 1648800000, 1648803600, 1648807200, 
    1648810800, 1648814400, 1648818000, 1648821600, 1648825200, 1648828800, 
    1648832400, 1648836000, 1648839600, 1648843200, 1648846800, 1648850400, 
    1648854000, 1648857600, 1648861200, 1648864800, 1648868400, 1648872000, 
    1648875600, 1648879200, 1648882800, 1648886400, 1648890000, 1648893600, 
    1648897200, 1648900800, 1648904400, 1648908000, 1648911600, 1648915200, 
    1648918800, 1648922400, 1648926000, 1648929600, 1648933200, 1648936800, 
    1648940400, 1648944000, 1648947600, 1648951200, 1648954800, 1648958400, 
    1648962000, 1648965600, 1648969200, 1648972800, 1648976400, 1648980000, 
    1648983600, 1648987200, 1648990800, 1648994400, 1648998000, 1649001600, 
    1649005200, 1649008800, 1649012400, 1649016000, 1649019600, 1649023200, 
    1649026800, 1649030400, 1649034000, 1649037600, 1649041200, 1649044800, 
    1649048400, 1649052000, 1649055600, 1649059200, 1649062800, 1649066400, 
    1649070000, 1649073600, 1649077200, 1649080800, 1649084400, 1649088000, 
    1649091600, 1649095200, 1649098800, 1649102400, 1649106000, 1649109600, 
    1649113200, 1649116800, 1649120400, 1649124000, 1649127600, 1649131200, 
    1649134800, 1649138400, 1649142000, 1649145600, 1649149200, 1649152800, 
    1649156400, 1649160000, 1649163600, 1649167200, 1649170800, 1649174400, 
    1649178000, 1649181600, 1649185200, 1649188800, 1649192400, 1649196000, 
    1649199600, 1649203200, 1649206800, 1649210400, 1649214000, 1649217600, 
    1649221200, 1649224800, 1649228400, 1649232000, 1649235600, 1649239200, 
    1649242800, 1649246400, 1649250000, 1649253600, 1649257200, 1649260800, 
    1649264400, 1649268000, 1649271600, 1649275200, 1649278800, 1649282400, 
    1649286000, 1649289600, 1649293200, 1649296800, 1649300400, 1649304000, 
    1649307600, 1649311200, 1649314800, 1649318400, 1649322000, 1649325600, 
    1649329200, 1649332800, 1649336400, 1649340000, 1649343600, 1649347200, 
    1649350800, 1649354400, 1649358000, 1649361600, 1649365200, 1649368800, 
    1649372400, 1649376000, 1649379600, 1649383200, 1649386800, 1649390400, 
    1649394000, 1649397600, 1649401200, 1649404800, 1649408400, 1649412000, 
    1649415600, 1649419200, 1649422800, 1649426400, 1649430000, 1649433600, 
    1649437200, 1649440800, 1649444400, 1649448000, 1649451600, 1649455200, 
    1649458800, 1649462400, 1649466000, 1649469600, 1649473200, 1649476800, 
    1649480400, 1649484000, 1649487600, 1649491200, 1649494800, 1649498400, 
    1649502000, 1649505600, 1649509200, 1649512800, 1649516400, 1649520000, 
    1649523600, 1649527200, 1649530800, 1649534400, 1649538000, 1649541600, 
    1649545200, 1649548800, 1649552400, 1649556000, 1649559600, 1649563200, 
    1649566800, 1649570400, 1649574000, 1649577600, 1649581200, 1649584800, 
    1649588400, 1649592000, 1649595600, 1649599200, 1649602800, 1649606400, 
    1649610000, 1649613600, 1649617200, 1649620800, 1649624400, 1649628000, 
    1649631600, 1649635200, 1649638800, 1649642400, 1649646000, 1649649600, 
    1649653200, 1649656800, 1649660400, 1649664000, 1649667600, 1649671200, 
    1649674800, 1649678400, 1649682000, 1649685600, 1649689200, 1649692800, 
    1649696400, 1649700000, 1649703600, 1649707200, 1649710800, 1649714400, 
    1649718000, 1649721600, 1649725200, 1649728800, 1649732400, 1649736000, 
    1649739600, 1649743200, 1649746800, 1649750400, 1649754000, 1649757600, 
    1649761200, 1649764800, 1649768400, 1649772000, 1649775600, 1649779200, 
    1649782800, 1649786400, 1649790000, 1649793600, 1649797200, 1649800800, 
    1649804400, 1649808000, 1649811600, 1649815200, 1649818800, 1649822400, 
    1649826000, 1649829600, 1649833200, 1649836800, 1649840400, 1649844000, 
    1649847600, 1649851200, 1649854800, 1649858400, 1649862000, 1649865600, 
    1649869200, 1649872800, 1649876400, 1649880000, 1649883600, 1649887200, 
    1649890800, 1649894400, 1649898000, 1649901600, 1649905200, 1649908800, 
    1649912400, 1649916000, 1649919600, 1649923200, 1649926800, 1649930400, 
    1649934000, 1649937600, 1649941200, 1649944800, 1649948400, 1649952000, 
    1649955600, 1649959200, 1649962800, 1649966400, 1649970000, 1649973600, 
    1649977200, 1649980800, 1649984400, 1649988000, 1649991600, 1649995200, 
    1649998800, 1650002400, 1650006000, 1650009600, 1650013200, 1650016800, 
    1650020400, 1650024000, 1650027600, 1650031200, 1650034800, 1650038400, 
    1650042000, 1650045600, 1650049200, 1650052800, 1650056400, 1650060000, 
    1650063600, 1650067200, 1650070800, 1650074400, 1650078000, 1650081600, 
    1650085200, 1650088800, 1650092400, 1650096000, 1650099600, 1650103200, 
    1650106800, 1650110400, 1650114000, 1650117600, 1650121200, 1650124800, 
    1650128400, 1650132000, 1650135600, 1650139200, 1650142800, 1650146400, 
    1650150000, 1650153600, 1650157200, 1650160800, 1650164400, 1650168000, 
    1650171600, 1650175200, 1650178800, 1650182400, 1650186000, 1650189600, 
    1650193200, 1650196800, 1650200400, 1650204000, 1650207600, 1650211200, 
    1650214800, 1650218400, 1650222000, 1650225600, 1650229200, 1650232800, 
    1650236400, 1650240000, 1650243600, 1650247200, 1650250800, 1650254400, 
    1650258000, 1650261600, 1650265200, 1650268800, 1650272400, 1650276000, 
    1650279600, 1650283200, 1650286800, 1650290400, 1650294000, 1650297600, 
    1650301200, 1650304800, 1650308400, 1650312000, 1650315600, 1650319200, 
    1650322800, 1650326400, 1650330000, 1650333600, 1650337200, 1650340800, 
    1650344400, 1650348000, 1650351600, 1650355200, 1650358800, 1650362400, 
    1650366000, 1650369600, 1650373200, 1650376800, 1650380400, 1650384000, 
    1650387600, 1650391200, 1650394800, 1650398400, 1650402000, 1650405600, 
    1650409200, 1650412800, 1650416400, 1650420000, 1650423600, 1650427200, 
    1650430800, 1650434400, 1650438000, 1650441600, 1650445200, 1650448800, 
    1650452400, 1650456000, 1650459600, 1650463200, 1650466800, 1650470400, 
    1650474000, 1650477600, 1650481200, 1650484800, 1650488400, 1650492000, 
    1650495600, 1650499200, 1650502800, 1650506400, 1650510000, 1650513600, 
    1650517200, 1650520800, 1650524400, 1650528000, 1650531600, 1650535200, 
    1650538800, 1650542400, 1650546000, 1650549600, 1650553200, 1650556800, 
    1650560400, 1650564000, 1650567600, 1650571200, 1650574800, 1650578400, 
    1650582000, 1650585600, 1650589200, 1650592800, 1650596400, 1650600000, 
    1650603600, 1650607200, 1650610800, 1650614400, 1650618000, 1650621600, 
    1650625200, 1650628800, 1650632400, 1650636000, 1650639600, 1650643200, 
    1650646800, 1650650400, 1650654000, 1650657600, 1650661200, 1650664800, 
    1650668400, 1650672000, 1650675600, 1650679200, 1650682800, 1650686400, 
    1650690000, 1650693600, 1650697200, 1650700800, 1650704400, 1650708000, 
    1650711600, 1650715200, 1650718800, 1650722400, 1650726000, 1650729600, 
    1650733200, 1650736800, 1650740400, 1650744000, 1650747600, 1650751200, 
    1650754800, 1650758400, 1650762000, 1650765600, 1650769200, 1650772800, 
    1650776400, 1650780000, 1650783600, 1650787200, 1650790800, 1650794400, 
    1650798000, 1650801600, 1650805200, 1650808800, 1650812400, 1650816000, 
    1650819600, 1650823200, 1650826800, 1650830400, 1650834000, 1650837600, 
    1650841200, 1650844800, 1650848400, 1650852000, 1650855600, 1650859200, 
    1650862800, 1650866400, 1650870000, 1650873600, 1650877200, 1650880800, 
    1650884400, 1650888000, 1650891600, 1650895200, 1650898800, 1650902400, 
    1650906000, 1650909600, 1650913200, 1650916800, 1650920400, 1650924000, 
    1650927600, 1650931200, 1650934800, 1650938400, 1650942000, 1650945600, 
    1650949200, 1650952800, 1650956400, 1650960000, 1650963600, 1650967200, 
    1650970800, 1650974400, 1650978000, 1650981600, 1650985200, 1650988800, 
    1650992400, 1650996000, 1650999600, 1651003200, 1651006800, 1651010400, 
    1651014000, 1651017600, 1651021200, 1651024800, 1651028400, 1651032000, 
    1651035600, 1651039200, 1651042800, 1651046400, 1651050000, 1651053600, 
    1651057200, 1651060800, 1651064400, 1651068000, 1651071600, 1651075200, 
    1651078800, 1651082400, 1651086000, 1651089600, 1651093200, 1651096800, 
    1651100400, 1651104000, 1651107600, 1651111200, 1651114800, 1651118400, 
    1651122000, 1651125600, 1651129200, 1651132800, 1651136400, 1651140000, 
    1651143600, 1651147200, 1651150800, 1651154400, 1651158000, 1651161600, 
    1651165200, 1651168800, 1651172400, 1651176000, 1651179600, 1651183200, 
    1651186800, 1651190400, 1651194000, 1651197600, 1651201200, 1651204800, 
    1651208400, 1651212000, 1651215600, 1651219200, 1651222800, 1651226400, 
    1651230000, 1651233600, 1651237200, 1651240800, 1651244400, 1651248000, 
    1651251600, 1651255200, 1651258800, 1651262400, 1651266000, 1651269600, 
    1651273200, 1651276800, 1651280400, 1651284000, 1651287600, 1651291200, 
    1651294800, 1651298400, 1651302000, 1651305600, 1651309200, 1651312800, 
    1651316400, 1651320000, 1651323600, 1651327200, 1651330800, 1651334400, 
    1651338000, 1651341600, 1651345200, 1651348800, 1651352400, 1651356000, 
    1651359600, 1651363200, 1651366800, 1651370400, 1651374000, 1651377600, 
    1651381200, 1651384800, 1651388400, 1651392000, 1651395600, 1651399200, 
    1651402800, 1651406400, 1651410000, 1651413600, 1651417200, 1651420800, 
    1651424400, 1651428000, 1651431600, 1651435200, 1651438800, 1651442400, 
    1651446000, 1651449600, 1651453200, 1651456800, 1651460400, 1651464000, 
    1651467600, 1651471200, 1651474800, 1651478400, 1651482000, 1651485600, 
    1651489200, 1651492800, 1651496400, 1651500000, 1651503600, 1651507200, 
    1651510800, 1651514400, 1651518000, 1651521600, 1651525200, 1651528800, 
    1651532400, 1651536000, 1651539600, 1651543200, 1651546800, 1651550400, 
    1651554000, 1651557600, 1651561200, 1651564800, 1651568400, 1651572000, 
    1651575600, 1651579200, 1651582800, 1651586400, 1651590000, 1651593600, 
    1651597200, 1651600800, 1651604400, 1651608000, 1651611600, 1651615200, 
    1651618800, 1651622400, 1651626000, 1651629600, 1651633200, 1651636800, 
    1651640400, 1651644000, 1651647600, 1651651200, 1651654800, 1651658400, 
    1651662000, 1651665600, 1651669200, 1651672800, 1651676400, 1651680000, 
    1651683600, 1651687200, 1651690800, 1651694400, 1651698000, 1651701600, 
    1651705200, 1651708800, 1651712400, 1651716000, 1651719600, 1651723200, 
    1651726800, 1651730400, 1651734000, 1651737600, 1651741200, 1651744800, 
    1651748400, 1651752000, 1651755600, 1651759200, 1651762800, 1651766400, 
    1651770000, 1651773600, 1651777200, 1651780800, 1651784400, 1651788000, 
    1651791600, 1651795200, 1651798800, 1651802400, 1651806000, 1651809600, 
    1651813200, 1651816800, 1651820400, 1651824000, 1651827600, 1651831200, 
    1651834800, 1651838400, 1651842000, 1651845600, 1651849200, 1651852800, 
    1651856400, 1651860000, 1651863600, 1651867200, 1651870800, 1651874400, 
    1651878000, 1651881600, 1651885200, 1651888800, 1651892400, 1651896000, 
    1651899600, 1651903200, 1651906800, 1651910400, 1651914000, 1651917600, 
    1651921200, 1651924800, 1651928400, 1651932000, 1651935600, 1651939200, 
    1651942800, 1651946400, 1651950000, 1651953600, 1651957200, 1651960800, 
    1651964400, 1651968000, 1651971600, 1651975200, 1651978800, 1651982400, 
    1651986000, 1651989600, 1651993200, 1651996800, 1652000400, 1652004000, 
    1652007600, 1652011200, 1652014800, 1652018400, 1652022000, 1652025600, 
    1652029200, 1652032800, 1652036400, 1652040000, 1652043600, 1652047200, 
    1652050800, 1652054400, 1652058000, 1652061600, 1652065200, 1652068800, 
    1652072400, 1652076000, 1652079600, 1652083200, 1652086800, 1652090400, 
    1652094000, 1652097600, 1652101200, 1652104800, 1652108400, 1652112000, 
    1652115600, 1652119200, 1652122800, 1652126400, 1652130000, 1652133600, 
    1652137200, 1652140800, 1652144400, 1652148000, 1652151600, 1652155200, 
    1652158800, 1652162400, 1652166000, 1652169600, 1652173200, 1652176800, 
    1652180400, 1652184000, 1652187600, 1652191200, 1652194800, 1652198400, 
    1652202000, 1652205600, 1652209200, 1652212800, 1652216400, 1652220000, 
    1652223600, 1652227200, 1652230800, 1652234400, 1652238000, 1652241600, 
    1652245200, 1652248800, 1652252400, 1652256000, 1652259600, 1652263200, 
    1652266800, 1652270400, 1652274000, 1652277600, 1652281200, 1652284800, 
    1652288400, 1652292000, 1652295600, 1652299200, 1652302800, 1652306400, 
    1652310000, 1652313600, 1652317200, 1652320800, 1652324400, 1652328000, 
    1652331600, 1652335200, 1652338800, 1652342400, 1652346000, 1652349600, 
    1652353200, 1652356800, 1652360400, 1652364000, 1652367600, 1652371200, 
    1652374800, 1652378400, 1652382000, 1652385600, 1652389200, 1652392800, 
    1652396400, 1652400000, 1652403600, 1652407200, 1652410800, 1652414400, 
    1652418000, 1652421600, 1652425200, 1652428800, 1652432400, 1652436000, 
    1652439600, 1652443200, 1652446800, 1652450400, 1652454000, 1652457600, 
    1652461200, 1652464800, 1652468400, 1652472000, 1652475600, 1652479200, 
    1652482800, 1652486400, 1652490000, 1652493600, 1652497200, 1652500800, 
    1652504400, 1652508000, 1652511600, 1652515200, 1652518800, 1652522400, 
    1652526000, 1652529600, 1652533200, 1652536800, 1652540400, 1652544000, 
    1652547600, 1652551200, 1652554800, 1652558400, 1652562000, 1652565600, 
    1652569200, 1652572800, 1652576400, 1652580000, 1652583600, 1652587200, 
    1652590800, 1652594400, 1652598000, 1652601600, 1652605200, 1652608800, 
    1652612400, 1652616000, 1652619600, 1652623200, 1652626800, 1652630400, 
    1652634000, 1652637600, 1652641200, 1652644800, 1652648400, 1652652000, 
    1652655600, 1652659200, 1652662800, 1652666400, 1652670000, 1652673600, 
    1652677200, 1652680800, 1652684400, 1652688000, 1652691600, 1652695200, 
    1652698800, 1652702400, 1652706000, 1652709600, 1652713200, 1652716800, 
    1652720400, 1652724000, 1652727600, 1652731200, 1652734800, 1652738400, 
    1652742000, 1652745600, 1652749200, 1652752800, 1652756400, 1652760000, 
    1652763600, 1652767200, 1652770800, 1652774400, 1652778000, 1652781600, 
    1652785200, 1652788800, 1652792400, 1652796000, 1652799600, 1652803200, 
    1652806800, 1652810400, 1652814000, 1652817600, 1652821200, 1652824800, 
    1652828400, 1652832000, 1652835600, 1652839200, 1652842800, 1652846400, 
    1652850000, 1652853600, 1652857200, 1652860800, 1652864400, 1652868000, 
    1652871600, 1652875200, 1652878800, 1652882400, 1652886000, 1652889600, 
    1652893200, 1652896800, 1652900400, 1652904000, 1652907600, 1652911200, 
    1652914800, 1652918400, 1652922000, 1652925600, 1652929200, 1652932800, 
    1652936400, 1652940000, 1652943600, 1652947200, 1652950800, 1652954400, 
    1652958000, 1652961600, 1652965200, 1652968800, 1652972400, 1652976000, 
    1652979600, 1652983200, 1652986800, 1652990400, 1652994000, 1652997600, 
    1653001200, 1653004800, 1653008400, 1653012000, 1653015600, 1653019200, 
    1653022800, 1653026400, 1653030000, 1653033600, 1653037200, 1653040800, 
    1653044400, 1653048000, 1653051600, 1653055200, 1653058800, 1653062400, 
    1653066000, 1653069600, 1653073200, 1653076800, 1653080400, 1653084000, 
    1653087600, 1653091200, 1653094800, 1653098400, 1653102000, 1653105600, 
    1653109200, 1653112800, 1653116400, 1653120000, 1653123600, 1653127200, 
    1653130800, 1653134400, 1653138000, 1653141600, 1653145200, 1653148800, 
    1653152400, 1653156000, 1653159600, 1653163200, 1653166800, 1653170400, 
    1653174000, 1653177600, 1653181200, 1653184800, 1653188400, 1653192000, 
    1653195600, 1653199200, 1653202800, 1653206400, 1653210000, 1653213600, 
    1653217200, 1653220800, 1653224400, 1653228000, 1653231600, 1653235200, 
    1653238800, 1653242400, 1653246000, 1653249600, 1653253200, 1653256800, 
    1653260400, 1653264000, 1653267600, 1653271200, 1653274800, 1653278400, 
    1653282000, 1653285600, 1653289200, 1653292800, 1653296400, 1653300000, 
    1653303600, 1653307200, 1653310800, 1653314400, 1653318000, 1653321600, 
    1653325200, 1653328800, 1653332400, 1653336000, 1653339600, 1653343200, 
    1653346800, 1653350400, 1653354000, 1653357600, 1653361200, 1653364800, 
    1653368400, 1653372000, 1653375600, 1653379200, 1653382800, 1653386400, 
    1653390000, 1653393600, 1653397200, 1653400800, 1653404400, 1653408000, 
    1653411600, 1653415200, 1653418800, 1653422400, 1653426000, 1653429600, 
    1653433200, 1653436800, 1653440400, 1653444000, 1653447600, 1653451200, 
    1653454800, 1653458400, 1653462000, 1653465600, 1653469200, 1653472800, 
    1653476400, 1653480000, 1653483600, 1653487200, 1653490800, 1653494400, 
    1653498000, 1653501600, 1653505200, 1653508800, 1653512400, 1653516000, 
    1653519600, 1653523200, 1653526800, 1653530400, 1653534000, 1653537600, 
    1653541200, 1653544800, 1653548400, 1653552000, 1653555600, 1653559200, 
    1653562800, 1653566400, 1653570000, 1653573600, 1653577200, 1653580800, 
    1653584400, 1653588000, 1653591600, 1653595200, 1653598800, 1653602400, 
    1653606000, 1653609600, 1653613200, 1653616800, 1653620400, 1653624000, 
    1653627600, 1653631200, 1653634800, 1653638400, 1653642000, 1653645600, 
    1653649200, 1653652800, 1653656400, 1653660000, 1653663600, 1653667200, 
    1653670800, 1653674400, 1653678000, 1653681600, 1653685200, 1653688800, 
    1653692400, 1653696000, 1653699600, 1653703200, 1653706800, 1653710400, 
    1653714000, 1653717600, 1653721200, 1653724800, 1653728400, 1653732000, 
    1653735600, 1653739200, 1653742800, 1653746400, 1653750000, 1653753600, 
    1653757200, 1653760800, 1653764400, 1653768000, 1653771600, 1653775200, 
    1653778800, 1653782400, 1653786000, 1653789600, 1653793200, 1653796800, 
    1653800400, 1653804000, 1653807600, 1653811200, 1653814800, 1653818400, 
    1653822000, 1653825600, 1653829200, 1653832800, 1653836400, 1653840000, 
    1653843600, 1653847200, 1653850800, 1653854400, 1653858000, 1653861600, 
    1653865200, 1653868800, 1653872400, 1653876000, 1653879600, 1653883200, 
    1653886800, 1653890400, 1653894000, 1653897600, 1653901200, 1653904800, 
    1653908400, 1653912000, 1653915600, 1653919200, 1653922800, 1653926400, 
    1653930000, 1653933600, 1653937200, 1653940800, 1653944400, 1653948000, 
    1653951600, 1653955200, 1653958800, 1653962400, 1653966000, 1653969600, 
    1653973200, 1653976800, 1653980400, 1653984000, 1653987600, 1653991200, 
    1653994800, 1653998400, 1654002000, 1654005600, 1654009200, 1654012800, 
    1654016400, 1654020000, 1654023600, 1654027200, 1654030800, 1654034400, 
    1654038000, 1654041600, 1654045200, 1654048800, 1654052400, 1654056000, 
    1654059600, 1654063200, 1654066800, 1654070400, 1654074000, 1654077600, 
    1654081200, 1654084800, 1654088400, 1654092000, 1654095600, 1654099200, 
    1654102800, 1654106400, 1654110000, 1654113600, 1654117200, 1654120800, 
    1654124400, 1654128000, 1654131600, 1654135200, 1654138800, 1654142400, 
    1654146000, 1654149600, 1654153200, 1654156800, 1654160400, 1654164000, 
    1654167600, 1654171200, 1654174800, 1654178400, 1654182000, 1654185600, 
    1654189200, 1654192800, 1654196400, 1654200000, 1654203600, 1654207200, 
    1654210800, 1654214400, 1654218000, 1654221600, 1654225200, 1654228800, 
    1654232400, 1654236000, 1654239600, 1654243200, 1654246800, 1654250400, 
    1654254000, 1654257600, 1654261200, 1654264800, 1654268400, 1654272000, 
    1654275600, 1654279200, 1654282800, 1654286400, 1654290000, 1654293600, 
    1654297200, 1654300800, 1654304400, 1654308000, 1654311600, 1654315200, 
    1654318800, 1654322400, 1654326000, 1654329600, 1654333200, 1654336800, 
    1654340400, 1654344000, 1654347600, 1654351200, 1654354800, 1654358400, 
    1654362000, 1654365600, 1654369200, 1654372800, 1654376400, 1654380000, 
    1654383600, 1654387200, 1654390800, 1654394400, 1654398000, 1654401600, 
    1654405200, 1654408800, 1654412400, 1654416000, 1654419600, 1654423200, 
    1654426800, 1654430400, 1654434000, 1654437600, 1654441200, 1654444800, 
    1654448400, 1654452000, 1654455600, 1654459200, 1654462800, 1654466400, 
    1654470000, 1654473600, 1654477200, 1654480800, 1654484400, 1654488000, 
    1654491600, 1654495200, 1654498800, 1654502400, 1654506000, 1654509600, 
    1654513200, 1654516800, 1654520400, 1654524000, 1654527600, 1654531200, 
    1654534800, 1654538400, 1654542000, 1654545600, 1654549200, 1654552800, 
    1654556400, 1654560000, 1654563600, 1654567200, 1654570800, 1654574400, 
    1654578000, 1654581600, 1654585200, 1654588800, 1654592400, 1654596000, 
    1654599600, 1654603200, 1654606800, 1654610400, 1654614000, 1654617600, 
    1654621200, 1654624800, 1654628400, 1654632000, 1654635600, 1654639200, 
    1654642800, 1654646400, 1654650000, 1654653600, 1654657200, 1654660800, 
    1654664400, 1654668000, 1654671600, 1654675200, 1654678800, 1654682400, 
    1654686000, 1654689600, 1654693200, 1654696800, 1654700400, 1654704000, 
    1654707600, 1654711200, 1654714800, 1654718400, 1654722000, 1654725600, 
    1654729200, 1654732800, 1654736400, 1654740000, 1654743600, 1654747200, 
    1654750800, 1654754400, 1654758000, 1654761600, 1654765200, 1654768800, 
    1654772400, 1654776000, 1654779600, 1654783200, 1654786800, 1654790400, 
    1654794000, 1654797600, 1654801200, 1654804800, 1654808400, 1654812000, 
    1654815600, 1654819200, 1654822800, 1654826400, 1654830000, 1654833600, 
    1654837200, 1654840800, 1654844400, 1654848000, 1654851600, 1654855200, 
    1654858800, 1654862400, 1654866000, 1654869600, 1654873200, 1654876800, 
    1654880400, 1654884000, 1654887600, 1654891200, 1654894800, 1654898400, 
    1654902000, 1654905600, 1654909200, 1654912800, 1654916400, 1654920000, 
    1654923600, 1654927200, 1654930800, 1654934400, 1654938000, 1654941600, 
    1654945200, 1654948800, 1654952400, 1654956000, 1654959600, 1654963200, 
    1654966800, 1654970400, 1654974000, 1654977600, 1654981200, 1654984800, 
    1654988400, 1654992000, 1654995600, 1654999200, 1655002800, 1655006400, 
    1655010000, 1655013600, 1655017200, 1655020800, 1655024400, 1655028000, 
    1655031600, 1655035200, 1655038800, 1655042400, 1655046000, 1655049600, 
    1655053200, 1655056800, 1655060400, 1655064000, 1655067600, 1655071200, 
    1655074800, 1655078400, 1655082000, 1655085600, 1655089200, 1655092800, 
    1655096400, 1655100000, 1655103600, 1655107200, 1655110800, 1655114400, 
    1655118000, 1655121600, 1655125200, 1655128800, 1655132400, 1655136000, 
    1655139600, 1655143200, 1655146800, 1655150400, 1655154000, 1655157600, 
    1655161200, 1655164800, 1655168400, 1655172000, 1655175600, 1655179200, 
    1655182800, 1655186400, 1655190000, 1655193600, 1655197200, 1655200800, 
    1655204400, 1655208000, 1655211600, 1655215200, 1655218800, 1655222400, 
    1655226000, 1655229600, 1655233200, 1655236800, 1655240400, 1655244000, 
    1655247600, 1655251200, 1655254800, 1655258400, 1655262000, 1655265600, 
    1655269200, 1655272800, 1655276400, 1655280000, 1655283600, 1655287200, 
    1655290800, 1655294400, 1655298000, 1655301600, 1655305200, 1655308800, 
    1655312400, 1655316000, 1655319600, 1655323200, 1655326800, 1655330400, 
    1655334000, 1655337600, 1655341200, 1655344800, 1655348400, 1655352000, 
    1655355600, 1655359200, 1655362800, 1655366400, 1655370000, 1655373600, 
    1655377200, 1655380800, 1655384400, 1655388000, 1655391600, 1655395200, 
    1655398800, 1655402400, 1655406000, 1655409600, 1655413200, 1655416800, 
    1655420400, 1655424000, 1655427600, 1655431200, 1655434800, 1655438400, 
    1655442000, 1655445600, 1655449200, 1655452800, 1655456400, 1655460000, 
    1655463600, 1655467200, 1655470800, 1655474400, 1655478000, 1655481600, 
    1655485200, 1655488800, 1655492400, 1655496000, 1655499600, 1655503200, 
    1655506800, 1655510400, 1655514000, 1655517600, 1655521200, 1655524800, 
    1655528400, 1655532000, 1655535600, 1655539200, 1655542800, 1655546400, 
    1655550000, 1655553600, 1655557200, 1655560800, 1655564400, 1655568000, 
    1655571600, 1655575200, 1655578800, 1655582400, 1655586000, 1655589600, 
    1655593200, 1655596800, 1655600400, 1655604000, 1655607600, 1655611200, 
    1655614800, 1655618400, 1655622000, 1655625600, 1655629200, 1655632800, 
    1655636400, 1655640000, 1655643600, 1655647200, 1655650800, 1655654400, 
    1655658000, 1655661600, 1655665200, 1655668800, 1655672400, 1655676000, 
    1655679600, 1655683200, 1655686800, 1655690400, 1655694000, 1655697600, 
    1655701200, 1655704800, 1655708400, 1655712000, 1655715600, 1655719200, 
    1655722800, 1655726400, 1655730000, 1655733600, 1655737200, 1655740800, 
    1655744400, 1655748000, 1655751600, 1655755200, 1655758800, 1655762400, 
    1655766000, 1655769600, 1655773200, 1655776800, 1655780400, 1655784000, 
    1655787600, 1655791200, 1655794800, 1655798400, 1655802000, 1655805600, 
    1655809200, 1655812800, 1655816400, 1655820000, 1655823600, 1655827200, 
    1655830800, 1655834400, 1655838000, 1655841600, 1655845200, 1655848800, 
    1655852400, 1655856000, 1655859600, 1655863200, 1655866800, 1655870400, 
    1655874000, 1655877600, 1655881200, 1655884800, 1655888400, 1655892000, 
    1655895600, 1655899200, 1655902800, 1655906400, 1655910000, 1655913600, 
    1655917200, 1655920800, 1655924400, 1655928000, 1655931600, 1655935200, 
    1655938800, 1655942400, 1655946000, 1655949600, 1655953200, 1655956800, 
    1655960400, 1655964000, 1655967600, 1655971200, 1655974800, 1655978400, 
    1655982000, 1655985600, 1655989200, 1655992800, 1655996400, 1656000000, 
    1656003600, 1656007200, 1656010800, 1656014400, 1656018000, 1656021600, 
    1656025200, 1656028800, 1656032400, 1656036000, 1656039600, 1656043200, 
    1656046800, 1656050400, 1656054000, 1656057600, 1656061200, 1656064800, 
    1656068400, 1656072000, 1656075600, 1656079200, 1656082800, 1656086400, 
    1656090000, 1656093600, 1656097200, 1656100800, 1656104400, 1656108000, 
    1656111600, 1656115200, 1656118800, 1656122400, 1656126000, 1656129600, 
    1656133200, 1656136800, 1656140400, 1656144000, 1656147600, 1656151200, 
    1656154800, 1656158400, 1656162000, 1656165600, 1656169200, 1656172800, 
    1656176400, 1656180000, 1656183600, 1656187200, 1656190800, 1656194400, 
    1656198000, 1656201600, 1656205200, 1656208800, 1656212400, 1656216000, 
    1656219600, 1656223200, 1656226800, 1656230400, 1656234000, 1656237600, 
    1656241200, 1656244800, 1656248400, 1656252000, 1656255600, 1656259200, 
    1656262800, 1656266400, 1656270000, 1656273600, 1656277200, 1656280800, 
    1656284400, 1656288000, 1656291600, 1656295200, 1656298800, 1656302400, 
    1656306000, 1656309600, 1656313200, 1656316800, 1656320400, 1656324000, 
    1656327600, 1656331200, 1656334800, 1656338400, 1656342000, 1656345600, 
    1656349200, 1656352800, 1656356400, 1656360000, 1656363600, 1656367200, 
    1656370800, 1656374400, 1656378000, 1656381600, 1656385200, 1656388800, 
    1656392400, 1656396000, 1656399600, 1656403200, 1656406800, 1656410400, 
    1656414000, 1656417600, 1656421200, 1656424800, 1656428400, 1656432000, 
    1656435600, 1656439200, 1656442800, 1656446400, 1656450000, 1656453600, 
    1656457200, 1656460800, 1656464400, 1656468000, 1656471600, 1656475200, 
    1656478800, 1656482400, 1656486000, 1656489600, 1656493200, 1656496800, 
    1656500400, 1656504000, 1656507600, 1656511200, 1656514800, 1656518400, 
    1656522000, 1656525600, 1656529200, 1656532800, 1656536400, 1656540000, 
    1656543600, 1656547200, 1656550800, 1656554400, 1656558000, 1656561600, 
    1656565200, 1656568800, 1656572400, 1656576000, 1656579600, 1656583200, 
    1656586800, 1656590400, 1656594000, 1656597600, 1656601200, 1656604800, 
    1656608400, 1656612000, 1656615600, 1656619200, 1656622800, 1656626400, 
    1656630000, 1656633600, 1656637200, 1656640800, 1656644400, 1656648000, 
    1656651600, 1656655200, 1656658800, 1656662400, 1656666000, 1656669600, 
    1656673200, 1656676800, 1656680400, 1656684000, 1656687600, 1656691200, 
    1656694800, 1656698400, 1656702000, 1656705600, 1656709200, 1656712800, 
    1656716400, 1656720000, 1656723600, 1656727200, 1656730800, 1656734400, 
    1656738000, 1656741600, 1656745200, 1656748800, 1656752400, 1656756000, 
    1656759600, 1656763200, 1656766800, 1656770400, 1656774000, 1656777600, 
    1656781200, 1656784800, 1656788400, 1656792000, 1656795600, 1656799200, 
    1656802800, 1656806400, 1656810000, 1656813600, 1656817200, 1656820800, 
    1656824400, 1656828000, 1656831600, 1656835200, 1656838800, 1656842400, 
    1656846000, 1656849600, 1656853200, 1656856800, 1656860400, 1656864000, 
    1656867600, 1656871200, 1656874800, 1656878400, 1656882000, 1656885600, 
    1656889200, 1656892800, 1656896400, 1656900000, 1656903600, 1656907200, 
    1656910800, 1656914400, 1656918000, 1656921600, 1656925200, 1656928800, 
    1656932400, 1656936000, 1656939600, 1656943200, 1656946800, 1656950400, 
    1656954000, 1656957600, 1656961200, 1656964800, 1656968400, 1656972000, 
    1656975600, 1656979200, 1656982800, 1656986400, 1656990000, 1656993600, 
    1656997200, 1657000800, 1657004400, 1657008000, 1657011600, 1657015200, 
    1657018800, 1657022400, 1657026000, 1657029600, 1657033200, 1657036800, 
    1657040400, 1657044000, 1657047600, 1657051200, 1657054800, 1657058400, 
    1657062000, 1657065600, 1657069200, 1657072800, 1657076400, 1657080000, 
    1657083600, 1657087200, 1657090800, 1657094400, 1657098000, 1657101600, 
    1657105200, 1657108800, 1657112400, 1657116000, 1657119600, 1657123200, 
    1657126800, 1657130400, 1657134000, 1657137600, 1657141200, 1657144800, 
    1657148400, 1657152000, 1657155600, 1657159200, 1657162800, 1657166400, 
    1657170000, 1657173600, 1657177200, 1657180800, 1657184400, 1657188000, 
    1657191600, 1657195200, 1657198800, 1657202400, 1657206000, 1657209600, 
    1657213200, 1657216800, 1657220400, 1657224000, 1657227600, 1657231200, 
    1657234800, 1657238400, 1657242000, 1657245600, 1657249200, 1657252800, 
    1657256400, 1657260000, 1657263600, 1657267200, 1657270800, 1657274400, 
    1657278000, 1657281600, 1657285200, 1657288800, 1657292400, 1657296000, 
    1657299600, 1657303200, 1657306800, 1657310400, 1657314000, 1657317600, 
    1657321200, 1657324800, 1657328400, 1657332000, 1657335600, 1657339200, 
    1657342800, 1657346400, 1657350000, 1657353600, 1657357200, 1657360800, 
    1657364400, 1657368000, 1657371600, 1657375200, 1657378800, 1657382400, 
    1657386000, 1657389600, 1657393200, 1657396800, 1657400400, 1657404000, 
    1657407600, 1657411200, 1657414800, 1657418400, 1657422000, 1657425600, 
    1657429200, 1657432800, 1657436400, 1657440000, 1657443600, 1657447200, 
    1657450800, 1657454400, 1657458000, 1657461600, 1657465200, 1657468800, 
    1657472400, 1657476000, 1657479600, 1657483200, 1657486800, 1657490400, 
    1657494000, 1657497600, 1657501200, 1657504800, 1657508400, 1657512000, 
    1657515600, 1657519200, 1657522800, 1657526400, 1657530000, 1657533600, 
    1657537200, 1657540800, 1657544400, 1657548000, 1657551600, 1657555200, 
    1657558800, 1657562400, 1657566000, 1657569600, 1657573200, 1657576800, 
    1657580400, 1657584000, 1657587600, 1657591200, 1657594800, 1657598400, 
    1657602000, 1657605600, 1657609200, 1657612800, 1657616400, 1657620000, 
    1657623600, 1657627200, 1657630800, 1657634400, 1657638000, 1657641600, 
    1657645200, 1657648800, 1657652400, 1657656000, 1657659600, 1657663200, 
    1657666800, 1657670400, 1657674000, 1657677600, 1657681200, 1657684800, 
    1657688400, 1657692000, 1657695600, 1657699200, 1657702800, 1657706400, 
    1657710000, 1657713600, 1657717200, 1657720800, 1657724400, 1657728000, 
    1657731600, 1657735200, 1657738800, 1657742400, 1657746000, 1657749600, 
    1657753200, 1657756800, 1657760400, 1657764000, 1657767600, 1657771200, 
    1657774800, 1657778400, 1657782000, 1657785600, 1657789200, 1657792800, 
    1657796400, 1657800000, 1657803600, 1657807200, 1657810800, 1657814400, 
    1657818000, 1657821600, 1657825200, 1657828800, 1657832400, 1657836000, 
    1657839600, 1657843200, 1657846800, 1657850400, 1657854000, 1657857600, 
    1657861200, 1657864800, 1657868400, 1657872000, 1657875600, 1657879200, 
    1657882800, 1657886400, 1657890000, 1657893600, 1657897200, 1657900800, 
    1657904400, 1657908000, 1657911600, 1657915200, 1657918800, 1657922400, 
    1657926000, 1657929600, 1657933200, 1657936800, 1657940400, 1657944000, 
    1657947600, 1657951200, 1657954800, 1657958400, 1657962000, 1657965600, 
    1657969200, 1657972800, 1657976400, 1657980000, 1657983600, 1657987200, 
    1657990800, 1657994400, 1657998000, 1658001600, 1658005200, 1658008800, 
    1658012400, 1658016000, 1658019600, 1658023200, 1658026800, 1658030400, 
    1658034000, 1658037600, 1658041200, 1658044800, 1658048400, 1658052000, 
    1658055600, 1658059200, 1658062800, 1658066400, 1658070000, 1658073600, 
    1658077200, 1658080800, 1658084400, 1658088000, 1658091600, 1658095200, 
    1658098800, 1658102400, 1658106000, 1658109600, 1658113200, 1658116800, 
    1658120400, 1658124000, 1658127600, 1658131200, 1658134800, 1658138400, 
    1658142000, 1658145600, 1658149200, 1658152800, 1658156400, 1658160000, 
    1658163600, 1658167200, 1658170800, 1658174400, 1658178000, 1658181600, 
    1658185200, 1658188800, 1658192400, 1658196000, 1658199600, 1658203200, 
    1658206800, 1658210400, 1658214000, 1658217600, 1658221200, 1658224800, 
    1658228400, 1658232000, 1658235600, 1658239200, 1658242800, 1658246400, 
    1658250000, 1658253600, 1658257200, 1658260800, 1658264400, 1658268000, 
    1658271600, 1658275200, 1658278800, 1658282400, 1658286000, 1658289600, 
    1658293200, 1658296800, 1658300400, 1658304000, 1658307600, 1658311200, 
    1658314800, 1658318400, 1658322000, 1658325600, 1658329200, 1658332800, 
    1658336400, 1658340000, 1658343600, 1658347200, 1658350800, 1658354400, 
    1658358000, 1658361600, 1658365200, 1658368800, 1658372400, 1658376000, 
    1658379600, 1658383200, 1658386800, 1658390400, 1658394000, 1658397600, 
    1658401200, 1658404800, 1658408400, 1658412000, 1658415600, 1658419200, 
    1658422800, 1658426400, 1658430000, 1658433600, 1658437200, 1658440800, 
    1658444400, 1658448000, 1658451600, 1658455200, 1658458800, 1658462400, 
    1658466000, 1658469600, 1658473200, 1658476800, 1658480400, 1658484000, 
    1658487600, 1658491200, 1658494800, 1658498400, 1658502000, 1658505600, 
    1658509200, 1658512800, 1658516400, 1658520000, 1658523600, 1658527200, 
    1658530800, 1658534400, 1658538000, 1658541600, 1658545200, 1658548800, 
    1658552400, 1658556000, 1658559600, 1658563200, 1658566800, 1658570400, 
    1658574000, 1658577600, 1658581200, 1658584800, 1658588400, 1658592000, 
    1658595600, 1658599200, 1658602800, 1658606400, 1658610000, 1658613600, 
    1658617200, 1658620800, 1658624400, 1658628000, 1658631600, 1658635200, 
    1658638800, 1658642400, 1658646000, 1658649600, 1658653200, 1658656800, 
    1658660400, 1658664000, 1658667600, 1658671200, 1658674800, 1658678400, 
    1658682000, 1658685600, 1658689200, 1658692800, 1658696400, 1658700000, 
    1658703600, 1658707200, 1658710800, 1658714400, 1658718000, 1658721600, 
    1658725200, 1658728800, 1658732400, 1658736000, 1658739600, 1658743200, 
    1658746800, 1658750400, 1658754000, 1658757600, 1658761200, 1658764800, 
    1658768400, 1658772000, 1658775600, 1658779200, 1658782800, 1658786400, 
    1658790000, 1658793600, 1658797200, 1658800800, 1658804400, 1658808000, 
    1658811600, 1658815200, 1658818800, 1658822400, 1658826000, 1658829600, 
    1658833200, 1658836800, 1658840400, 1658844000, 1658847600, 1658851200, 
    1658854800, 1658858400, 1658862000, 1658865600, 1658869200, 1658872800, 
    1658876400, 1658880000, 1658883600, 1658887200, 1658890800, 1658894400, 
    1658898000, 1658901600, 1658905200, 1658908800, 1658912400, 1658916000, 
    1658919600, 1658923200, 1658926800, 1658930400, 1658934000, 1658937600, 
    1658941200, 1658944800, 1658948400, 1658952000, 1658955600, 1658959200, 
    1658962800, 1658966400, 1658970000, 1658973600, 1658977200, 1658980800, 
    1658984400, 1658988000, 1658991600, 1658995200, 1658998800, 1659002400, 
    1659006000, 1659009600, 1659013200, 1659016800, 1659020400, 1659024000, 
    1659027600, 1659031200, 1659034800, 1659038400, 1659042000, 1659045600, 
    1659049200, 1659052800, 1659056400, 1659060000, 1659063600, 1659067200, 
    1659070800, 1659074400, 1659078000, 1659081600, 1659085200, 1659088800, 
    1659092400, 1659096000, 1659099600, 1659103200, 1659106800, 1659110400, 
    1659114000, 1659117600, 1659121200, 1659124800, 1659128400, 1659132000, 
    1659135600, 1659139200, 1659142800, 1659146400, 1659150000, 1659153600, 
    1659157200, 1659160800, 1659164400, 1659168000, 1659171600, 1659175200, 
    1659178800, 1659182400, 1659186000, 1659189600, 1659193200, 1659196800, 
    1659200400, 1659204000, 1659207600, 1659211200, 1659214800, 1659218400, 
    1659222000, 1659225600, 1659229200, 1659232800, 1659236400, 1659240000, 
    1659243600, 1659247200, 1659250800, 1659254400, 1659258000, 1659261600, 
    1659265200, 1659268800, 1659272400, 1659276000, 1659279600, 1659283200, 
    1659286800, 1659290400, 1659294000, 1659297600, 1659301200, 1659304800, 
    1659308400, 1659312000, 1659315600, 1659319200, 1659322800, 1659326400, 
    1659330000, 1659333600, 1659337200, 1659340800, 1659344400, 1659348000, 
    1659351600, 1659355200, 1659358800, 1659362400, 1659366000, 1659369600, 
    1659373200, 1659376800, 1659380400, 1659384000, 1659387600, 1659391200, 
    1659394800, 1659398400, 1659402000, 1659405600, 1659409200, 1659412800, 
    1659416400, 1659420000, 1659423600, 1659427200, 1659430800, 1659434400, 
    1659438000, 1659441600, 1659445200, 1659448800, 1659452400, 1659456000, 
    1659459600, 1659463200, 1659466800, 1659470400, 1659474000, 1659477600, 
    1659481200, 1659484800, 1659488400, 1659492000, 1659495600, 1659499200, 
    1659502800, 1659506400, 1659510000, 1659513600, 1659517200, 1659520800, 
    1659524400, 1659528000, 1659531600, 1659535200, 1659538800, 1659542400, 
    1659546000, 1659549600, 1659553200, 1659556800, 1659560400, 1659564000, 
    1659567600, 1659571200, 1659574800, 1659578400, 1659582000, 1659585600, 
    1659589200, 1659592800, 1659596400, 1659600000, 1659603600, 1659607200, 
    1659610800, 1659614400, 1659618000, 1659621600, 1659625200, 1659628800, 
    1659632400, 1659636000, 1659639600, 1659643200, 1659646800, 1659650400, 
    1659654000, 1659657600, 1659661200, 1659664800, 1659668400, 1659672000, 
    1659675600, 1659679200, 1659682800, 1659686400, 1659690000, 1659693600, 
    1659697200, 1659700800, 1659704400, 1659708000, 1659711600, 1659715200, 
    1659718800, 1659722400, 1659726000, 1659729600, 1659733200, 1659736800, 
    1659740400, 1659744000, 1659747600, 1659751200, 1659754800, 1659758400, 
    1659762000, 1659765600, 1659769200, 1659772800, 1659776400, 1659780000, 
    1659783600, 1659787200, 1659790800, 1659794400, 1659798000, 1659801600, 
    1659805200, 1659808800, 1659812400, 1659816000, 1659819600, 1659823200, 
    1659826800, 1659830400, 1659834000, 1659837600, 1659841200, 1659844800, 
    1659848400, 1659852000, 1659855600, 1659859200, 1659862800, 1659866400, 
    1659870000, 1659873600, 1659877200, 1659880800, 1659884400, 1659888000, 
    1659891600, 1659895200, 1659898800, 1659902400, 1659906000, 1659909600, 
    1659913200, 1659916800, 1659920400, 1659924000, 1659927600, 1659931200, 
    1659934800, 1659938400, 1659942000, 1659945600, 1659949200, 1659952800, 
    1659956400, 1659960000, 1659963600, 1659967200, 1659970800, 1659974400, 
    1659978000, 1659981600, 1659985200, 1659988800, 1659992400, 1659996000, 
    1659999600, 1660003200, 1660006800, 1660010400, 1660014000, 1660017600, 
    1660021200, 1660024800, 1660028400, 1660032000, 1660035600, 1660039200, 
    1660042800, 1660046400, 1660050000, 1660053600, 1660057200, 1660060800, 
    1660064400, 1660068000, 1660071600, 1660075200, 1660078800, 1660082400, 
    1660086000, 1660089600, 1660093200, 1660096800, 1660100400, 1660104000, 
    1660107600, 1660111200, 1660114800, 1660118400, 1660122000, 1660125600, 
    1660129200, 1660132800, 1660136400, 1660140000, 1660143600, 1660147200, 
    1660150800, 1660154400, 1660158000, 1660161600, 1660165200, 1660168800, 
    1660172400, 1660176000, 1660179600, 1660183200, 1660186800, 1660190400, 
    1660194000, 1660197600, 1660201200, 1660204800, 1660208400, 1660212000, 
    1660215600, 1660219200, 1660222800, 1660226400, 1660230000, 1660233600, 
    1660237200, 1660240800, 1660244400, 1660248000, 1660251600, 1660255200, 
    1660258800, 1660262400, 1660266000, 1660269600, 1660273200, 1660276800, 
    1660280400, 1660284000, 1660287600, 1660291200, 1660294800, 1660298400, 
    1660302000, 1660305600, 1660309200, 1660312800, 1660316400, 1660320000, 
    1660323600, 1660327200, 1660330800, 1660334400, 1660338000, 1660341600, 
    1660345200, 1660348800, 1660352400, 1660356000, 1660359600, 1660363200, 
    1660366800, 1660370400, 1660374000, 1660377600, 1660381200, 1660384800, 
    1660388400, 1660392000, 1660395600, 1660399200, 1660402800, 1660406400, 
    1660410000, 1660413600, 1660417200, 1660420800, 1660424400, 1660428000, 
    1660431600, 1660435200, 1660438800, 1660442400, 1660446000, 1660449600, 
    1660453200, 1660456800, 1660460400, 1660464000, 1660467600, 1660471200, 
    1660474800, 1660478400, 1660482000, 1660485600, 1660489200, 1660492800, 
    1660496400, 1660500000, 1660503600, 1660507200, 1660510800, 1660514400, 
    1660518000, 1660521600, 1660525200, 1660528800, 1660532400, 1660536000, 
    1660539600, 1660543200, 1660546800, 1660550400, 1660554000, 1660557600, 
    1660561200, 1660564800, 1660568400, 1660572000, 1660575600, 1660579200, 
    1660582800, 1660586400, 1660590000, 1660593600, 1660597200, 1660600800, 
    1660604400, 1660608000, 1660611600, 1660615200, 1660618800, 1660622400, 
    1660626000, 1660629600, 1660633200, 1660636800, 1660640400, 1660644000, 
    1660647600, 1660651200, 1660654800, 1660658400, 1660662000, 1660665600, 
    1660669200, 1660672800, 1660676400, 1660680000, 1660683600, 1660687200, 
    1660690800, 1660694400, 1660698000, 1660701600, 1660705200, 1660708800, 
    1660712400, 1660716000, 1660719600, 1660723200, 1660726800, 1660730400, 
    1660734000, 1660737600, 1660741200, 1660744800, 1660748400, 1660752000, 
    1660755600, 1660759200, 1660762800, 1660766400, 1660770000, 1660773600, 
    1660777200, 1660780800, 1660784400, 1660788000, 1660791600, 1660795200, 
    1660798800, 1660802400, 1660806000, 1660809600, 1660813200, 1660816800, 
    1660820400, 1660824000, 1660827600, 1660831200, 1660834800, 1660838400, 
    1660842000, 1660845600, 1660849200, 1660852800, 1660856400, 1660860000, 
    1660863600, 1660867200, 1660870800, 1660874400, 1660878000, 1660881600, 
    1660885200, 1660888800, 1660892400, 1660896000, 1660899600, 1660903200, 
    1660906800, 1660910400, 1660914000, 1660917600, 1660921200, 1660924800, 
    1660928400, 1660932000, 1660935600, 1660939200, 1660942800, 1660946400, 
    1660950000, 1660953600, 1660957200, 1660960800, 1660964400, 1660968000, 
    1660971600, 1660975200, 1660978800, 1660982400, 1660986000, 1660989600, 
    1660993200, 1660996800, 1661000400, 1661004000, 1661007600, 1661011200, 
    1661014800, 1661018400, 1661022000, 1661025600, 1661029200, 1661032800, 
    1661036400, 1661040000, 1661043600, 1661047200, 1661050800, 1661054400, 
    1661058000, 1661061600, 1661065200, 1661068800, 1661072400, 1661076000, 
    1661079600, 1661083200, 1661086800, 1661090400, 1661094000, 1661097600, 
    1661101200, 1661104800, 1661108400, 1661112000, 1661115600, 1661119200, 
    1661122800, 1661126400, 1661130000, 1661133600, 1661137200, 1661140800, 
    1661144400, 1661148000, 1661151600, 1661155200, 1661158800, 1661162400, 
    1661166000, 1661169600, 1661173200, 1661176800, 1661180400, 1661184000, 
    1661187600, 1661191200, 1661194800, 1661198400, 1661202000, 1661205600, 
    1661209200, 1661212800, 1661216400, 1661220000, 1661223600, 1661227200, 
    1661230800, 1661234400, 1661238000, 1661241600, 1661245200, 1661248800, 
    1661252400, 1661256000, 1661259600, 1661263200, 1661266800, 1661270400, 
    1661274000, 1661277600, 1661281200, 1661284800, 1661288400, 1661292000, 
    1661295600, 1661299200, 1661302800, 1661306400, 1661310000, 1661313600, 
    1661317200, 1661320800, 1661324400, 1661328000, 1661331600, 1661335200, 
    1661338800, 1661342400, 1661346000, 1661349600, 1661353200, 1661356800, 
    1661360400, 1661364000, 1661367600, 1661371200, 1661374800, 1661378400, 
    1661382000, 1661385600, 1661389200, 1661392800, 1661396400, 1661400000, 
    1661403600, 1661407200, 1661410800, 1661414400, 1661418000, 1661421600, 
    1661425200, 1661428800, 1661432400, 1661436000, 1661439600, 1661443200, 
    1661446800, 1661450400, 1661454000, 1661457600, 1661461200, 1661464800, 
    1661468400, 1661472000, 1661475600, 1661479200, 1661482800, 1661486400, 
    1661490000, 1661493600, 1661497200, 1661500800, 1661504400, 1661508000, 
    1661511600, 1661515200, 1661518800, 1661522400, 1661526000, 1661529600, 
    1661533200, 1661536800, 1661540400, 1661544000, 1661547600, 1661551200, 
    1661554800, 1661558400, 1661562000, 1661565600, 1661569200, 1661572800, 
    1661576400, 1661580000, 1661583600, 1661587200, 1661590800, 1661594400, 
    1661598000, 1661601600, 1661605200, 1661608800, 1661612400, 1661616000, 
    1661619600, 1661623200, 1661626800, 1661630400, 1661634000, 1661637600, 
    1661641200, 1661644800, 1661648400, 1661652000, 1661655600, 1661659200, 
    1661662800, 1661666400, 1661670000, 1661673600, 1661677200, 1661680800, 
    1661684400, 1661688000, 1661691600, 1661695200, 1661698800, 1661702400, 
    1661706000, 1661709600, 1661713200, 1661716800, 1661720400, 1661724000, 
    1661727600, 1661731200, 1661734800, 1661738400, 1661742000, 1661745600, 
    1661749200, 1661752800, 1661756400, 1661760000, 1661763600, 1661767200, 
    1661770800, 1661774400, 1661778000, 1661781600, 1661785200, 1661788800, 
    1661792400, 1661796000, 1661799600, 1661803200, 1661806800, 1661810400, 
    1661814000, 1661817600, 1661821200, 1661824800, 1661828400, 1661832000, 
    1661835600, 1661839200, 1661842800, 1661846400, 1661850000, 1661853600, 
    1661857200, 1661860800, 1661864400, 1661868000, 1661871600, 1661875200, 
    1661878800, 1661882400, 1661886000, 1661889600, 1661893200, 1661896800, 
    1661900400, 1661904000, 1661907600, 1661911200, 1661914800, 1661918400, 
    1661922000, 1661925600, 1661929200, 1661932800, 1661936400, 1661940000, 
    1661943600, 1661947200, 1661950800, 1661954400, 1661958000, 1661961600, 
    1661965200, 1661968800, 1661972400, 1661976000, 1661979600, 1661983200, 
    1661986800, 1661990400, 1661994000, 1661997600, 1662001200, 1662004800, 
    1662008400, 1662012000, 1662015600, 1662019200, 1662022800, 1662026400, 
    1662030000, 1662033600, 1662037200, 1662040800, 1662044400, 1662048000, 
    1662051600, 1662055200, 1662058800, 1662062400, 1662066000, 1662069600, 
    1662073200, 1662076800, 1662080400, 1662084000, 1662087600, 1662091200, 
    1662094800, 1662098400, 1662102000, 1662105600, 1662109200, 1662112800, 
    1662116400, 1662120000, 1662123600, 1662127200, 1662130800, 1662134400, 
    1662138000, 1662141600, 1662145200, 1662148800, 1662152400, 1662156000, 
    1662159600, 1662163200, 1662166800, 1662170400, 1662174000, 1662177600, 
    1662181200, 1662184800, 1662188400, 1662192000, 1662195600, 1662199200, 
    1662202800, 1662206400, 1662210000, 1662213600, 1662217200, 1662220800, 
    1662224400, 1662228000, 1662231600, 1662235200, 1662238800, 1662242400, 
    1662246000, 1662249600, 1662253200, 1662256800, 1662260400, 1662264000, 
    1662267600, 1662271200, 1662274800, 1662278400, 1662282000, 1662285600, 
    1662289200, 1662292800, 1662296400, 1662300000, 1662303600, 1662307200, 
    1662310800, 1662314400, 1662318000, 1662321600, 1662325200, 1662328800, 
    1662332400, 1662336000, 1662339600, 1662343200, 1662346800, 1662350400, 
    1662354000, 1662357600, 1662361200, 1662364800, 1662368400, 1662372000, 
    1662375600, 1662379200, 1662382800, 1662386400, 1662390000, 1662393600, 
    1662397200, 1662400800, 1662404400, 1662408000, 1662411600, 1662415200, 
    1662418800, 1662422400, 1662426000, 1662429600, 1662433200, 1662436800, 
    1662440400, 1662444000, 1662447600, 1662451200, 1662454800, 1662458400, 
    1662462000, 1662465600, 1662469200, 1662472800, 1662476400, 1662480000, 
    1662483600, 1662487200, 1662490800, 1662494400, 1662498000, 1662501600, 
    1662505200, 1662508800, 1662512400, 1662516000, 1662519600, 1662523200, 
    1662526800, 1662530400, 1662534000, 1662537600, 1662541200, 1662544800, 
    1662548400, 1662552000, 1662555600, 1662559200, 1662562800, 1662566400, 
    1662570000, 1662573600, 1662577200, 1662580800, 1662584400, 1662588000, 
    1662591600, 1662595200, 1662598800, 1662602400, 1662606000, 1662609600, 
    1662613200, 1662616800, 1662620400, 1662624000, 1662627600, 1662631200, 
    1662634800, 1662638400, 1662642000, 1662645600, 1662649200, 1662652800, 
    1662656400, 1662660000, 1662663600, 1662667200, 1662670800, 1662674400, 
    1662678000, 1662681600, 1662685200, 1662688800, 1662692400, 1662696000, 
    1662699600, 1662703200, 1662706800, 1662710400, 1662714000, 1662717600, 
    1662721200, 1662724800, 1662728400, 1662732000, 1662735600, 1662739200, 
    1662742800, 1662746400, 1662750000, 1662753600, 1662757200, 1662760800, 
    1662764400, 1662768000, 1662771600, 1662775200, 1662778800, 1662782400, 
    1662786000, 1662789600, 1662793200, 1662796800, 1662800400, 1662804000, 
    1662807600, 1662811200, 1662814800, 1662818400, 1662822000, 1662825600, 
    1662829200, 1662832800, 1662836400, 1662840000, 1662843600, 1662847200, 
    1662850800, 1662854400, 1662858000, 1662861600, 1662865200, 1662868800, 
    1662872400, 1662876000, 1662879600, 1662883200, 1662886800, 1662890400, 
    1662894000, 1662897600, 1662901200, 1662904800, 1662908400, 1662912000, 
    1662915600, 1662919200, 1662922800, 1662926400, 1662930000, 1662933600, 
    1662937200, 1662940800, 1662944400, 1662948000, 1662951600, 1662955200, 
    1662958800, 1662962400, 1662966000, 1662969600, 1662973200, 1662976800, 
    1662980400, 1662984000, 1662987600, 1662991200, 1662994800, 1662998400, 
    1663002000, 1663005600, 1663009200, 1663012800, 1663016400, 1663020000, 
    1663023600, 1663027200, 1663030800, 1663034400, 1663038000, 1663041600, 
    1663045200, 1663048800, 1663052400, 1663056000, 1663059600, 1663063200, 
    1663066800, 1663070400, 1663074000, 1663077600, 1663081200, 1663084800, 
    1663088400, 1663092000, 1663095600, 1663099200, 1663102800, 1663106400, 
    1663110000, 1663113600, 1663117200, 1663120800, 1663124400, 1663128000, 
    1663131600, 1663135200, 1663138800, 1663142400, 1663146000, 1663149600, 
    1663153200, 1663156800, 1663160400, 1663164000, 1663167600, 1663171200, 
    1663174800, 1663178400, 1663182000, 1663185600, 1663189200, 1663192800, 
    1663196400, 1663200000, 1663203600, 1663207200, 1663210800, 1663214400, 
    1663218000, 1663221600, 1663225200, 1663228800, 1663232400, 1663236000, 
    1663239600, 1663243200, 1663246800, 1663250400, 1663254000, 1663257600, 
    1663261200, 1663264800, 1663268400, 1663272000, 1663275600, 1663279200, 
    1663282800, 1663286400, 1663290000, 1663293600, 1663297200, 1663300800, 
    1663304400, 1663308000, 1663311600, 1663315200, 1663318800, 1663322400, 
    1663326000, 1663329600, 1663333200, 1663336800, 1663340400, 1663344000, 
    1663347600, 1663351200, 1663354800, 1663358400, 1663362000, 1663365600, 
    1663369200, 1663372800, 1663376400, 1663380000, 1663383600, 1663387200, 
    1663390800, 1663394400, 1663398000, 1663401600, 1663405200, 1663408800, 
    1663412400, 1663416000, 1663419600, 1663423200, 1663426800, 1663430400, 
    1663434000, 1663437600, 1663441200, 1663444800, 1663448400, 1663452000, 
    1663455600, 1663459200, 1663462800, 1663466400, 1663470000, 1663473600, 
    1663477200, 1663480800, 1663484400, 1663488000, 1663491600, 1663495200, 
    1663498800, 1663502400, 1663506000, 1663509600, 1663513200, 1663516800, 
    1663520400, 1663524000, 1663527600, 1663531200, 1663534800, 1663538400, 
    1663542000, 1663545600, 1663549200, 1663552800, 1663556400, 1663560000, 
    1663563600, 1663567200, 1663570800, 1663574400, 1663578000, 1663581600, 
    1663585200, 1663588800, 1663592400, 1663596000, 1663599600, 1663603200, 
    1663606800, 1663610400, 1663614000, 1663617600, 1663621200, 1663624800, 
    1663628400, 1663632000, 1663635600, 1663639200, 1663642800, 1663646400, 
    1663650000, 1663653600, 1663657200, 1663660800, 1663664400, 1663668000, 
    1663671600, 1663675200, 1663678800, 1663682400, 1663686000, 1663689600, 
    1663693200, 1663696800, 1663700400, 1663704000, 1663707600, 1663711200, 
    1663714800, 1663718400, 1663722000, 1663725600, 1663729200, 1663732800, 
    1663736400, 1663740000, 1663743600, 1663747200, 1663750800, 1663754400, 
    1663758000, 1663761600, 1663765200, 1663768800, 1663772400, 1663776000, 
    1663779600, 1663783200, 1663786800, 1663790400, 1663794000, 1663797600, 
    1663801200, 1663804800, 1663808400, 1663812000, 1663815600, 1663819200, 
    1663822800, 1663826400, 1663830000, 1663833600, 1663837200, 1663840800, 
    1663844400, 1663848000, 1663851600, 1663855200, 1663858800, 1663862400, 
    1663866000, 1663869600, 1663873200, 1663876800, 1663880400, 1663884000, 
    1663887600, 1663891200, 1663894800, 1663898400, 1663902000, 1663905600, 
    1663909200, 1663912800, 1663916400, 1663920000, 1663923600, 1663927200, 
    1663930800, 1663934400, 1663938000, 1663941600, 1663945200, 1663948800, 
    1663952400, 1663956000, 1663959600, 1663963200, 1663966800, 1663970400, 
    1663974000, 1663977600, 1663981200, 1663984800, 1663988400, 1663992000, 
    1663995600, 1663999200, 1664002800, 1664006400, 1664010000, 1664013600, 
    1664017200, 1664020800, 1664024400, 1664028000, 1664031600, 1664035200, 
    1664038800, 1664042400, 1664046000, 1664049600, 1664053200, 1664056800, 
    1664060400, 1664064000, 1664067600, 1664071200, 1664074800, 1664078400, 
    1664082000, 1664085600, 1664089200, 1664092800, 1664096400, 1664100000, 
    1664103600, 1664107200, 1664110800, 1664114400, 1664118000, 1664121600, 
    1664125200, 1664128800, 1664132400, 1664136000, 1664139600, 1664143200, 
    1664146800, 1664150400, 1664154000, 1664157600, 1664161200, 1664164800, 
    1664168400, 1664172000, 1664175600, 1664179200, 1664182800, 1664186400, 
    1664190000, 1664193600, 1664197200, 1664200800, 1664204400, 1664208000, 
    1664211600, 1664215200, 1664218800, 1664222400, 1664226000, 1664229600, 
    1664233200, 1664236800, 1664240400, 1664244000, 1664247600, 1664251200, 
    1664254800, 1664258400, 1664262000, 1664265600, 1664269200, 1664272800, 
    1664276400, 1664280000, 1664283600, 1664287200, 1664290800, 1664294400, 
    1664298000, 1664301600, 1664305200, 1664308800, 1664312400, 1664316000, 
    1664319600, 1664323200, 1664326800, 1664330400, 1664334000, 1664337600, 
    1664341200, 1664344800, 1664348400, 1664352000, 1664355600, 1664359200, 
    1664362800, 1664366400, 1664370000, 1664373600, 1664377200, 1664380800, 
    1664384400, 1664388000, 1664391600, 1664395200, 1664398800, 1664402400, 
    1664406000, 1664409600, 1664413200, 1664416800, 1664420400, 1664424000, 
    1664427600, 1664431200, 1664434800, 1664438400, 1664442000, 1664445600, 
    1664449200, 1664452800, 1664456400, 1664460000, 1664463600, 1664467200, 
    1664470800, 1664474400, 1664478000, 1664481600, 1664485200, 1664488800, 
    1664492400, 1664496000, 1664499600, 1664503200, 1664506800, 1664510400, 
    1664514000, 1664517600, 1664521200, 1664524800, 1664528400, 1664532000, 
    1664535600, 1664539200, 1664542800, 1664546400, 1664550000, 1664553600, 
    1664557200, 1664560800, 1664564400, 1664568000, 1664571600, 1664575200, 
    1664578800, 1664582400, 1664586000, 1664589600, 1664593200, 1664596800, 
    1664600400, 1664604000, 1664607600, 1664611200, 1664614800, 1664618400, 
    1664622000, 1664625600, 1664629200, 1664632800, 1664636400, 1664640000, 
    1664643600, 1664647200, 1664650800, 1664654400, 1664658000, 1664661600, 
    1664665200, 1664668800, 1664672400, 1664676000, 1664679600, 1664683200, 
    1664686800, 1664690400, 1664694000, 1664697600, 1664701200, 1664704800, 
    1664708400, 1664712000, 1664715600, 1664719200, 1664722800, 1664726400, 
    1664730000, 1664733600, 1664737200, 1664740800, 1664744400, 1664748000, 
    1664751600, 1664755200, 1664758800, 1664762400, 1664766000, 1664769600, 
    1664773200, 1664776800, 1664780400, 1664784000, 1664787600, 1664791200, 
    1664794800, 1664798400, 1664802000, 1664805600, 1664809200, 1664812800, 
    1664816400, 1664820000, 1664823600, 1664827200, 1664830800, 1664834400, 
    1664838000, 1664841600, 1664845200, 1664848800, 1664852400, 1664856000, 
    1664859600, 1664863200, 1664866800, 1664870400, 1664874000, 1664877600, 
    1664881200, 1664884800, 1664888400, 1664892000, 1664895600, 1664899200, 
    1664902800, 1664906400, 1664910000, 1664913600, 1664917200, 1664920800, 
    1664924400, 1664928000, 1664931600, 1664935200, 1664938800, 1664942400, 
    1664946000, 1664949600, 1664953200, 1664956800, 1664960400, 1664964000, 
    1664967600, 1664971200, 1664974800, 1664978400, 1664982000, 1664985600, 
    1664989200, 1664992800, 1664996400, 1665000000, 1665003600, 1665007200, 
    1665010800, 1665014400, 1665018000, 1665021600, 1665025200, 1665028800, 
    1665032400, 1665036000, 1665039600, 1665043200, 1665046800, 1665050400, 
    1665054000, 1665057600, 1665061200, 1665064800, 1665068400, 1665072000, 
    1665075600, 1665079200, 1665082800, 1665086400, 1665090000, 1665093600, 
    1665097200, 1665100800, 1665104400, 1665108000, 1665111600, 1665115200, 
    1665118800, 1665122400, 1665126000, 1665129600, 1665133200, 1665136800, 
    1665140400, 1665144000, 1665147600, 1665151200, 1665154800, 1665158400, 
    1665162000, 1665165600, 1665169200, 1665172800, 1665176400, 1665180000, 
    1665183600, 1665187200, 1665190800, 1665194400, 1665198000, 1665201600, 
    1665205200, 1665208800, 1665212400, 1665216000, 1665219600, 1665223200, 
    1665226800, 1665230400, 1665234000, 1665237600, 1665241200, 1665244800, 
    1665248400, 1665252000, 1665255600, 1665259200, 1665262800, 1665266400, 
    1665270000, 1665273600, 1665277200, 1665280800, 1665284400, 1665288000, 
    1665291600, 1665295200, 1665298800, 1665302400, 1665306000, 1665309600, 
    1665313200, 1665316800, 1665320400, 1665324000, 1665327600, 1665331200, 
    1665334800, 1665338400, 1665342000, 1665345600, 1665349200, 1665352800, 
    1665356400, 1665360000, 1665363600, 1665367200, 1665370800, 1665374400, 
    1665378000, 1665381600, 1665385200, 1665388800, 1665392400, 1665396000, 
    1665399600, 1665403200, 1665406800, 1665410400, 1665414000, 1665417600, 
    1665421200, 1665424800, 1665428400, 1665432000, 1665435600, 1665439200, 
    1665442800, 1665446400, 1665450000, 1665453600, 1665457200, 1665460800, 
    1665464400, 1665468000, 1665471600, 1665475200, 1665478800, 1665482400, 
    1665486000, 1665489600, 1665493200, 1665496800, 1665500400, 1665504000, 
    1665507600, 1665511200, 1665514800, 1665518400, 1665522000, 1665525600, 
    1665529200, 1665532800, 1665536400, 1665540000, 1665543600, 1665547200, 
    1665550800, 1665554400, 1665558000, 1665561600, 1665565200, 1665568800, 
    1665572400, 1665576000, 1665579600, 1665583200, 1665586800, 1665590400, 
    1665594000, 1665597600, 1665601200, 1665604800, 1665608400, 1665612000, 
    1665615600, 1665619200, 1665622800, 1665626400, 1665630000, 1665633600, 
    1665637200, 1665640800, 1665644400, 1665648000, 1665651600, 1665655200, 
    1665658800, 1665662400, 1665666000, 1665669600, 1665673200, 1665676800, 
    1665680400, 1665684000, 1665687600, 1665691200, 1665694800, 1665698400, 
    1665702000, 1665705600, 1665709200, 1665712800, 1665716400, 1665720000, 
    1665723600, 1665727200, 1665730800, 1665734400, 1665738000, 1665741600, 
    1665745200, 1665748800, 1665752400, 1665756000, 1665759600, 1665763200, 
    1665766800, 1665770400, 1665774000, 1665777600, 1665781200, 1665784800, 
    1665788400, 1665792000, 1665795600, 1665799200, 1665802800, 1665806400, 
    1665810000, 1665813600, 1665817200, 1665820800, 1665824400, 1665828000, 
    1665831600, 1665835200, 1665838800, 1665842400, 1665846000, 1665849600, 
    1665853200, 1665856800, 1665860400, 1665864000, 1665867600, 1665871200, 
    1665874800, 1665878400, 1665882000, 1665885600, 1665889200, 1665892800, 
    1665896400, 1665900000, 1665903600, 1665907200, 1665910800, 1665914400, 
    1665918000, 1665921600, 1665925200, 1665928800, 1665932400, 1665936000, 
    1665939600, 1665943200, 1665946800, 1665950400, 1665954000, 1665957600, 
    1665961200, 1665964800, 1665968400, 1665972000, 1665975600, 1665979200, 
    1665982800, 1665986400, 1665990000, 1665993600, 1665997200, 1666000800, 
    1666004400, 1666008000, 1666011600, 1666015200, 1666018800, 1666022400, 
    1666026000, 1666029600, 1666033200, 1666036800, 1666040400, 1666044000, 
    1666047600, 1666051200, 1666054800, 1666058400, 1666062000, 1666065600, 
    1666069200, 1666072800, 1666076400, 1666080000, 1666083600, 1666087200, 
    1666090800, 1666094400, 1666098000, 1666101600, 1666105200, 1666108800, 
    1666112400, 1666116000, 1666119600, 1666123200, 1666126800, 1666130400, 
    1666134000, 1666137600, 1666141200, 1666144800, 1666148400, 1666152000, 
    1666155600, 1666159200, 1666162800, 1666166400, 1666170000, 1666173600, 
    1666177200, 1666180800, 1666184400, 1666188000, 1666191600, 1666195200, 
    1666198800, 1666202400, 1666206000, 1666209600, 1666213200, 1666216800, 
    1666220400, 1666224000, 1666227600, 1666231200, 1666234800, 1666238400, 
    1666242000, 1666245600, 1666249200, 1666252800, 1666256400, 1666260000, 
    1666263600, 1666267200, 1666270800, 1666274400, 1666278000, 1666281600, 
    1666285200, 1666288800, 1666292400, 1666296000, 1666299600, 1666303200, 
    1666306800, 1666310400, 1666314000, 1666317600, 1666321200, 1666324800, 
    1666328400, 1666332000, 1666335600, 1666339200, 1666342800, 1666346400, 
    1666350000, 1666353600, 1666357200, 1666360800, 1666364400, 1666368000, 
    1666371600, 1666375200, 1666378800, 1666382400, 1666386000, 1666389600, 
    1666393200, 1666396800, 1666400400, 1666404000, 1666407600, 1666411200, 
    1666414800, 1666418400, 1666422000, 1666425600, 1666429200, 1666432800, 
    1666436400, 1666440000, 1666443600, 1666447200, 1666450800, 1666454400, 
    1666458000, 1666461600, 1666465200, 1666468800, 1666472400, 1666476000, 
    1666479600, 1666483200, 1666486800, 1666490400, 1666494000, 1666497600, 
    1666501200, 1666504800, 1666508400, 1666512000, 1666515600, 1666519200, 
    1666522800, 1666526400, 1666530000, 1666533600, 1666537200, 1666540800, 
    1666544400, 1666548000, 1666551600, 1666555200, 1666558800, 1666562400, 
    1666566000, 1666569600, 1666573200, 1666576800, 1666580400, 1666584000, 
    1666587600, 1666591200, 1666594800, 1666598400, 1666602000, 1666605600, 
    1666609200, 1666612800, 1666616400, 1666620000, 1666623600, 1666627200, 
    1666630800, 1666634400, 1666638000, 1666641600, 1666645200, 1666648800, 
    1666652400, 1666656000, 1666659600, 1666663200, 1666666800, 1666670400, 
    1666674000, 1666677600, 1666681200, 1666684800, 1666688400, 1666692000, 
    1666695600, 1666699200, 1666702800, 1666706400, 1666710000, 1666713600, 
    1666717200, 1666720800, 1666724400, 1666728000, 1666731600, 1666735200, 
    1666738800, 1666742400, 1666746000, 1666749600, 1666753200, 1666756800, 
    1666760400, 1666764000, 1666767600, 1666771200, 1666774800, 1666778400, 
    1666782000, 1666785600, 1666789200, 1666792800, 1666796400, 1666800000, 
    1666803600, 1666807200, 1666810800, 1666814400, 1666818000, 1666821600, 
    1666825200, 1666828800, 1666832400, 1666836000, 1666839600, 1666843200, 
    1666846800, 1666850400, 1666854000, 1666857600, 1666861200, 1666864800, 
    1666868400, 1666872000, 1666875600, 1666879200, 1666882800, 1666886400, 
    1666890000, 1666893600, 1666897200, 1666900800, 1666904400, 1666908000, 
    1666911600, 1666915200, 1666918800, 1666922400, 1666926000, 1666929600, 
    1666933200, 1666936800, 1666940400, 1666944000, 1666947600, 1666951200, 
    1666954800, 1666958400, 1666962000, 1666965600, 1666969200, 1666972800, 
    1666976400, 1666980000, 1666983600, 1666987200, 1666990800, 1666994400, 
    1666998000, 1667001600, 1667005200, 1667008800, 1667012400, 1667016000, 
    1667019600, 1667023200, 1667026800, 1667030400, 1667034000, 1667037600, 
    1667041200, 1667044800, 1667048400, 1667052000, 1667055600, 1667059200, 
    1667062800, 1667066400, 1667070000, 1667073600, 1667077200, 1667080800, 
    1667084400, 1667088000, 1667091600, 1667095200, 1667098800, 1667102400, 
    1667106000, 1667109600, 1667113200, 1667116800, 1667120400, 1667124000, 
    1667127600, 1667131200, 1667134800, 1667138400, 1667142000, 1667145600, 
    1667149200, 1667152800, 1667156400, 1667160000, 1667163600, 1667167200, 
    1667170800, 1667174400, 1667178000, 1667181600, 1667185200, 1667188800, 
    1667192400, 1667196000, 1667199600, 1667203200, 1667206800, 1667210400, 
    1667214000, 1667217600, 1667221200, 1667224800, 1667228400, 1667232000, 
    1667235600, 1667239200, 1667242800, 1667246400, 1667250000, 1667253600, 
    1667257200, 1667260800, 1667264400, 1667268000, 1667271600, 1667275200, 
    1667278800, 1667282400, 1667286000, 1667289600, 1667293200, 1667296800, 
    1667300400, 1667304000, 1667307600, 1667311200, 1667314800, 1667318400, 
    1667322000, 1667325600, 1667329200, 1667332800, 1667336400, 1667340000, 
    1667343600, 1667347200, 1667350800, 1667354400, 1667358000, 1667361600, 
    1667365200, 1667368800, 1667372400, 1667376000, 1667379600, 1667383200, 
    1667386800, 1667390400, 1667394000, 1667397600, 1667401200, 1667404800, 
    1667408400, 1667412000, 1667415600, 1667419200, 1667422800, 1667426400, 
    1667430000, 1667433600, 1667437200, 1667440800, 1667444400, 1667448000, 
    1667451600, 1667455200, 1667458800, 1667462400, 1667466000, 1667469600, 
    1667473200, 1667476800, 1667480400, 1667484000, 1667487600, 1667491200, 
    1667494800, 1667498400, 1667502000, 1667505600, 1667509200, 1667512800, 
    1667516400, 1667520000, 1667523600, 1667527200, 1667530800, 1667534400, 
    1667538000, 1667541600, 1667545200, 1667548800, 1667552400, 1667556000, 
    1667559600, 1667563200, 1667566800, 1667570400, 1667574000, 1667577600, 
    1667581200, 1667584800, 1667588400, 1667592000, 1667595600, 1667599200, 
    1667602800, 1667606400, 1667610000, 1667613600, 1667617200, 1667620800, 
    1667624400, 1667628000, 1667631600, 1667635200, 1667638800, 1667642400, 
    1667646000, 1667649600, 1667653200, 1667656800, 1667660400, 1667664000, 
    1667667600, 1667671200, 1667674800, 1667678400, 1667682000, 1667685600, 
    1667689200, 1667692800, 1667696400, 1667700000, 1667703600, 1667707200, 
    1667710800, 1667714400, 1667718000, 1667721600, 1667725200, 1667728800, 
    1667732400, 1667736000, 1667739600, 1667743200, 1667746800, 1667750400, 
    1667754000, 1667757600, 1667761200, 1667764800, 1667768400, 1667772000, 
    1667775600, 1667779200, 1667782800, 1667786400, 1667790000, 1667793600, 
    1667797200, 1667800800, 1667804400, 1667808000, 1667811600, 1667815200, 
    1667818800, 1667822400, 1667826000, 1667829600, 1667833200, 1667836800, 
    1667840400, 1667844000, 1667847600, 1667851200, 1667854800, 1667858400, 
    1667862000, 1667865600, 1667869200, 1667872800, 1667876400, 1667880000, 
    1667883600, 1667887200, 1667890800, 1667894400, 1667898000, 1667901600, 
    1667905200, 1667908800, 1667912400, 1667916000, 1667919600, 1667923200, 
    1667926800, 1667930400, 1667934000, 1667937600, 1667941200, 1667944800, 
    1667948400, 1667952000, 1667955600, 1667959200, 1667962800, 1667966400, 
    1667970000, 1667973600, 1667977200, 1667980800, 1667984400, 1667988000, 
    1667991600, 1667995200, 1667998800, 1668002400, 1668006000, 1668009600, 
    1668013200, 1668016800, 1668020400, 1668024000, 1668027600, 1668031200, 
    1668034800, 1668038400, 1668042000, 1668045600, 1668049200, 1668052800, 
    1668056400, 1668060000, 1668063600, 1668067200, 1668070800, 1668074400, 
    1668078000, 1668081600, 1668085200, 1668088800, 1668092400, 1668096000, 
    1668099600, 1668103200, 1668106800, 1668110400, 1668114000, 1668117600, 
    1668121200, 1668124800, 1668128400, 1668132000, 1668135600, 1668139200, 
    1668142800, 1668146400, 1668150000, 1668153600, 1668157200, 1668160800, 
    1668164400, 1668168000, 1668171600, 1668175200, 1668178800, 1668182400, 
    1668186000, 1668189600, 1668193200, 1668196800, 1668200400, 1668204000, 
    1668207600, 1668211200, 1668214800, 1668218400, 1668222000, 1668225600, 
    1668229200, 1668232800, 1668236400, 1668240000, 1668243600, 1668247200, 
    1668250800, 1668254400, 1668258000, 1668261600, 1668265200, 1668268800, 
    1668272400, 1668276000, 1668279600, 1668283200, 1668286800, 1668290400, 
    1668294000, 1668297600, 1668301200, 1668304800, 1668308400, 1668312000, 
    1668315600, 1668319200, 1668322800, 1668326400, 1668330000, 1668333600, 
    1668337200, 1668340800, 1668344400, 1668348000, 1668351600, 1668355200, 
    1668358800, 1668362400, 1668366000, 1668369600, 1668373200, 1668376800, 
    1668380400, 1668384000, 1668387600, 1668391200, 1668394800, 1668398400, 
    1668402000, 1668405600, 1668409200, 1668412800, 1668416400, 1668420000, 
    1668423600, 1668427200, 1668430800, 1668434400, 1668438000, 1668441600, 
    1668445200, 1668448800, 1668452400, 1668456000, 1668459600, 1668463200, 
    1668466800, 1668470400, 1668474000, 1668477600, 1668481200, 1668484800, 
    1668488400, 1668492000, 1668495600, 1668499200, 1668502800, 1668506400, 
    1668510000, 1668513600, 1668517200, 1668520800, 1668524400, 1668528000, 
    1668531600, 1668535200, 1668538800, 1668542400, 1668546000, 1668549600, 
    1668553200, 1668556800, 1668560400, 1668564000, 1668567600, 1668571200, 
    1668574800, 1668578400, 1668582000, 1668585600, 1668589200, 1668592800, 
    1668596400, 1668600000, 1668603600, 1668607200, 1668610800, 1668614400, 
    1668618000, 1668621600, 1668625200, 1668628800, 1668632400, 1668636000, 
    1668639600, 1668643200, 1668646800, 1668650400, 1668654000, 1668657600, 
    1668661200, 1668664800, 1668668400, 1668672000, 1668675600, 1668679200, 
    1668682800, 1668686400, 1668690000, 1668693600, 1668697200, 1668700800, 
    1668704400, 1668708000, 1668711600, 1668715200, 1668718800, 1668722400, 
    1668726000, 1668729600, 1668733200, 1668736800, 1668740400, 1668744000, 
    1668747600, 1668751200, 1668754800, 1668758400, 1668762000, 1668765600, 
    1668769200, 1668772800, 1668776400, 1668780000, 1668783600, 1668787200, 
    1668790800, 1668794400, 1668798000, 1668801600, 1668805200, 1668808800, 
    1668812400, 1668816000, 1668819600, 1668823200, 1668826800, 1668830400, 
    1668834000, 1668837600, 1668841200, 1668844800, 1668848400, 1668852000, 
    1668855600, 1668859200, 1668862800, 1668866400, 1668870000, 1668873600, 
    1668877200, 1668880800, 1668884400, 1668888000, 1668891600, 1668895200, 
    1668898800, 1668902400, 1668906000, 1668909600, 1668913200, 1668916800, 
    1668920400, 1668924000, 1668927600, 1668931200, 1668934800, 1668938400, 
    1668942000, 1668945600, 1668949200, 1668952800, 1668956400, 1668960000, 
    1668963600, 1668967200, 1668970800, 1668974400, 1668978000, 1668981600, 
    1668985200, 1668988800, 1668992400, 1668996000, 1668999600, 1669003200, 
    1669006800, 1669010400, 1669014000, 1669017600, 1669021200, 1669024800, 
    1669028400, 1669032000, 1669035600, 1669039200, 1669042800, 1669046400, 
    1669050000, 1669053600, 1669057200, 1669060800, 1669064400, 1669068000, 
    1669071600, 1669075200, 1669078800, 1669082400, 1669086000, 1669089600, 
    1669093200, 1669096800, 1669100400, 1669104000, 1669107600, 1669111200, 
    1669114800, 1669118400, 1669122000, 1669125600, 1669129200, 1669132800, 
    1669136400, 1669140000, 1669143600, 1669147200, 1669150800, 1669154400, 
    1669158000, 1669161600, 1669165200, 1669168800, 1669172400, 1669176000, 
    1669179600, 1669183200, 1669186800, 1669190400, 1669194000, 1669197600, 
    1669201200, 1669204800, 1669208400, 1669212000, 1669215600, 1669219200, 
    1669222800, 1669226400, 1669230000, 1669233600, 1669237200, 1669240800, 
    1669244400, 1669248000, 1669251600, 1669255200, 1669258800, 1669262400, 
    1669266000, 1669269600, 1669273200, 1669276800, 1669280400, 1669284000, 
    1669287600, 1669291200, 1669294800, 1669298400, 1669302000, 1669305600, 
    1669309200, 1669312800, 1669316400, 1669320000, 1669323600, 1669327200, 
    1669330800, 1669334400, 1669338000, 1669341600, 1669345200, 1669348800, 
    1669352400, 1669356000, 1669359600, 1669363200, 1669366800, 1669370400, 
    1669374000, 1669377600, 1669381200, 1669384800, 1669388400, 1669392000, 
    1669395600, 1669399200, 1669402800, 1669406400, 1669410000, 1669413600, 
    1669417200, 1669420800, 1669424400, 1669428000, 1669431600, 1669435200, 
    1669438800, 1669442400, 1669446000, 1669449600, 1669453200, 1669456800, 
    1669460400, 1669464000, 1669467600, 1669471200, 1669474800, 1669478400, 
    1669482000, 1669485600, 1669489200, 1669492800, 1669496400, 1669500000, 
    1669503600, 1669507200, 1669510800, 1669514400, 1669518000, 1669521600, 
    1669525200, 1669528800, 1669532400, 1669536000, 1669539600, 1669543200, 
    1669546800, 1669550400, 1669554000, 1669557600, 1669561200, 1669564800, 
    1669568400, 1669572000, 1669575600, 1669579200, 1669582800, 1669586400, 
    1669590000, 1669593600, 1669597200, 1669600800, 1669604400, 1669608000, 
    1669611600, 1669615200, 1669618800, 1669622400, 1669626000, 1669629600, 
    1669633200, 1669636800, 1669640400, 1669644000, 1669647600, 1669651200, 
    1669654800, 1669658400, 1669662000, 1669665600, 1669669200, 1669672800, 
    1669676400, 1669680000, 1669683600, 1669687200, 1669690800, 1669694400, 
    1669698000, 1669701600, 1669705200, 1669708800, 1669712400, 1669716000, 
    1669719600, 1669723200, 1669726800, 1669730400, 1669734000, 1669737600, 
    1669741200, 1669744800, 1669748400, 1669752000, 1669755600, 1669759200, 
    1669762800, 1669766400, 1669770000, 1669773600, 1669777200, 1669780800, 
    1669784400, 1669788000, 1669791600, 1669795200, 1669798800, 1669802400, 
    1669806000, 1669809600, 1669813200, 1669816800, 1669820400, 1669824000, 
    1669827600, 1669831200, 1669834800, 1669838400, 1669842000, 1669845600, 
    1669849200, 1669852800, 1669856400, 1669860000, 1669863600, 1669867200, 
    1669870800, 1669874400, 1669878000, 1669881600, 1669885200, 1669888800, 
    1669892400, 1669896000, 1669899600, 1669903200, 1669906800, 1669910400, 
    1669914000, 1669917600, 1669921200, 1669924800, 1669928400, 1669932000, 
    1669935600, 1669939200, 1669942800, 1669946400, 1669950000, 1669953600, 
    1669957200, 1669960800, 1669964400, 1669968000, 1669971600, 1669975200, 
    1669978800, 1669982400, 1669986000, 1669989600, 1669993200, 1669996800, 
    1670000400, 1670004000, 1670007600, 1670011200, 1670014800, 1670018400, 
    1670022000, 1670025600, 1670029200, 1670032800, 1670036400, 1670040000, 
    1670043600, 1670047200, 1670050800, 1670054400, 1670058000, 1670061600, 
    1670065200, 1670068800, 1670072400, 1670076000, 1670079600, 1670083200, 
    1670086800, 1670090400, 1670094000, 1670097600, 1670101200, 1670104800, 
    1670108400, 1670112000, 1670115600, 1670119200, 1670122800, 1670126400, 
    1670130000, 1670133600, 1670137200, 1670140800, 1670144400, 1670148000, 
    1670151600, 1670155200, 1670158800, 1670162400, 1670166000, 1670169600, 
    1670173200, 1670176800, 1670180400, 1670184000, 1670187600, 1670191200, 
    1670194800, 1670198400, 1670202000, 1670205600, 1670209200, 1670212800, 
    1670216400, 1670220000, 1670223600, 1670227200, 1670230800, 1670234400, 
    1670238000, 1670241600, 1670245200, 1670248800, 1670252400, 1670256000, 
    1670259600, 1670263200, 1670266800, 1670270400, 1670274000, 1670277600, 
    1670281200, 1670284800, 1670288400, 1670292000, 1670295600, 1670299200, 
    1670302800, 1670306400, 1670310000, 1670313600, 1670317200, 1670320800, 
    1670324400, 1670328000, 1670331600, 1670335200, 1670338800, 1670342400, 
    1670346000, 1670349600, 1670353200, 1670356800, 1670360400, 1670364000, 
    1670367600, 1670371200, 1670374800, 1670378400, 1670382000, 1670385600, 
    1670389200, 1670392800, 1670396400, 1670400000, 1670403600, 1670407200, 
    1670410800, 1670414400, 1670418000, 1670421600, 1670425200, 1670428800, 
    1670432400, 1670436000, 1670439600, 1670443200, 1670446800, 1670450400, 
    1670454000, 1670457600, 1670461200, 1670464800, 1670468400, 1670472000, 
    1670475600, 1670479200, 1670482800, 1670486400, 1670490000, 1670493600, 
    1670497200, 1670500800, 1670504400, 1670508000, 1670511600, 1670515200, 
    1670518800, 1670522400, 1670526000, 1670529600, 1670533200, 1670536800, 
    1670540400, 1670544000, 1670547600, 1670551200, 1670554800, 1670558400, 
    1670562000, 1670565600, 1670569200, 1670572800, 1670576400, 1670580000, 
    1670583600, 1670587200, 1670590800, 1670594400, 1670598000, 1670601600, 
    1670605200, 1670608800, 1670612400, 1670616000, 1670619600, 1670623200, 
    1670626800, 1670630400, 1670634000, 1670637600, 1670641200, 1670644800, 
    1670648400, 1670652000, 1670655600, 1670659200, 1670662800, 1670666400, 
    1670670000, 1670673600, 1670677200, 1670680800, 1670684400, 1670688000, 
    1670691600, 1670695200, 1670698800, 1670702400, 1670706000, 1670709600, 
    1670713200, 1670716800, 1670720400, 1670724000, 1670727600, 1670731200, 
    1670734800, 1670738400, 1670742000, 1670745600, 1670749200, 1670752800, 
    1670756400, 1670760000, 1670763600, 1670767200, 1670770800, 1670774400, 
    1670778000, 1670781600, 1670785200, 1670788800, 1670792400, 1670796000, 
    1670799600, 1670803200, 1670806800, 1670810400, 1670814000, 1670817600, 
    1670821200, 1670824800, 1670828400, 1670832000, 1670835600, 1670839200, 
    1670842800, 1670846400, 1670850000, 1670853600, 1670857200, 1670860800, 
    1670864400, 1670868000, 1670871600, 1670875200, 1670878800, 1670882400, 
    1670886000, 1670889600, 1670893200, 1670896800, 1670900400, 1670904000, 
    1670907600, 1670911200, 1670914800, 1670918400, 1670922000, 1670925600, 
    1670929200, 1670932800, 1670936400, 1670940000, 1670943600, 1670947200, 
    1670950800, 1670954400, 1670958000, 1670961600, 1670965200, 1670968800, 
    1670972400, 1670976000, 1670979600, 1670983200, 1670986800, 1670990400, 
    1670994000, 1670997600, 1671001200, 1671004800, 1671008400, 1671012000, 
    1671015600, 1671019200, 1671022800, 1671026400, 1671030000, 1671033600, 
    1671037200, 1671040800, 1671044400, 1671048000, 1671051600, 1671055200, 
    1671058800, 1671062400, 1671066000, 1671069600, 1671073200, 1671076800, 
    1671080400, 1671084000, 1671087600, 1671091200, 1671094800, 1671098400, 
    1671102000, 1671105600, 1671109200, 1671112800, 1671116400, 1671120000, 
    1671123600, 1671127200, 1671130800, 1671134400, 1671138000, 1671141600, 
    1671145200, 1671148800, 1671152400, 1671156000, 1671159600, 1671163200, 
    1671166800, 1671170400, 1671174000, 1671177600, 1671181200, 1671184800, 
    1671188400, 1671192000, 1671195600, 1671199200, 1671202800, 1671206400, 
    1671210000, 1671213600, 1671217200, 1671220800, 1671224400, 1671228000, 
    1671231600, 1671235200, 1671238800, 1671242400, 1671246000, 1671249600, 
    1671253200, 1671256800, 1671260400, 1671264000, 1671267600, 1671271200, 
    1671274800, 1671278400, 1671282000, 1671285600, 1671289200, 1671292800, 
    1671296400, 1671300000, 1671303600, 1671307200, 1671310800, 1671314400, 
    1671318000, 1671321600, 1671325200, 1671328800, 1671332400, 1671336000, 
    1671339600, 1671343200, 1671346800, 1671350400, 1671354000, 1671357600, 
    1671361200, 1671364800, 1671368400, 1671372000, 1671375600, 1671379200, 
    1671382800, 1671386400, 1671390000, 1671393600, 1671397200, 1671400800, 
    1671404400, 1671408000, 1671411600, 1671415200, 1671418800, 1671422400, 
    1671426000, 1671429600, 1671433200, 1671436800, 1671440400, 1671444000, 
    1671447600, 1671451200, 1671454800, 1671458400, 1671462000, 1671465600, 
    1671469200, 1671472800, 1671476400, 1671480000, 1671483600, 1671487200, 
    1671490800, 1671494400, 1671498000, 1671501600, 1671505200, 1671508800, 
    1671512400, 1671516000, 1671519600, 1671523200, 1671526800, 1671530400, 
    1671534000, 1671537600, 1671541200, 1671544800, 1671548400, 1671552000, 
    1671555600, 1671559200, 1671562800, 1671566400, 1671570000, 1671573600, 
    1671577200, 1671580800, 1671584400, 1671588000, 1671591600, 1671595200, 
    1671598800, 1671602400, 1671606000, 1671609600, 1671613200, 1671616800, 
    1671620400, 1671624000, 1671627600, 1671631200, 1671634800, 1671638400, 
    1671642000, 1671645600, 1671649200, 1671652800, 1671656400, 1671660000, 
    1671663600, 1671667200, 1671670800, 1671674400, 1671678000, 1671681600, 
    1671685200, 1671688800, 1671692400, 1671696000, 1671699600, 1671703200, 
    1671706800, 1671710400, 1671714000, 1671717600, 1671721200, 1671724800, 
    1671728400, 1671732000, 1671735600, 1671739200, 1671742800, 1671746400, 
    1671750000, 1671753600, 1671757200, 1671760800, 1671764400, 1671768000, 
    1671771600, 1671775200, 1671778800, 1671782400, 1671786000, 1671789600, 
    1671793200, 1671796800, 1671800400, 1671804000, 1671807600, 1671811200, 
    1671814800, 1671818400, 1671822000, 1671825600, 1671829200, 1671832800, 
    1671836400, 1671840000, 1671843600, 1671847200, 1671850800, 1671854400, 
    1671858000, 1671861600, 1671865200, 1671868800, 1671872400, 1671876000, 
    1671879600, 1671883200, 1671886800, 1671890400, 1671894000, 1671897600, 
    1671901200, 1671904800, 1671908400, 1671912000, 1671915600, 1671919200, 
    1671922800, 1671926400, 1671930000, 1671933600, 1671937200, 1671940800, 
    1671944400, 1671948000, 1671951600, 1671955200, 1671958800, 1671962400, 
    1671966000, 1671969600, 1671973200, 1671976800, 1671980400, 1671984000, 
    1671987600, 1671991200, 1671994800, 1671998400, 1672002000, 1672005600, 
    1672009200, 1672012800, 1672016400, 1672020000, 1672023600, 1672027200, 
    1672030800, 1672034400, 1672038000, 1672041600, 1672045200, 1672048800, 
    1672052400, 1672056000, 1672059600, 1672063200, 1672066800, 1672070400, 
    1672074000, 1672077600, 1672081200, 1672084800, 1672088400, 1672092000, 
    1672095600, 1672099200, 1672102800, 1672106400, 1672110000, 1672113600, 
    1672117200, 1672120800, 1672124400, 1672128000, 1672131600, 1672135200, 
    1672138800, 1672142400, 1672146000, 1672149600, 1672153200, 1672156800, 
    1672160400, 1672164000, 1672167600, 1672171200, 1672174800, 1672178400, 
    1672182000, 1672185600, 1672189200, 1672192800, 1672196400, 1672200000, 
    1672203600, 1672207200, 1672210800, 1672214400, 1672218000, 1672221600, 
    1672225200, 1672228800, 1672232400, 1672236000, 1672239600, 1672243200, 
    1672246800, 1672250400, 1672254000, 1672257600, 1672261200, 1672264800, 
    1672268400, 1672272000, 1672275600, 1672279200, 1672282800, 1672286400, 
    1672290000, 1672293600, 1672297200, 1672300800, 1672304400, 1672308000, 
    1672311600, 1672315200, 1672318800, 1672322400, 1672326000, 1672329600, 
    1672333200, 1672336800, 1672340400, 1672344000, 1672347600, 1672351200, 
    1672354800, 1672358400, 1672362000, 1672365600, 1672369200, 1672372800, 
    1672376400, 1672380000, 1672383600, 1672387200, 1672390800, 1672394400, 
    1672398000, 1672401600, 1672405200, 1672408800, 1672412400, 1672416000, 
    1672419600, 1672423200, 1672426800, 1672430400, 1672434000, 1672437600, 
    1672441200, 1672444800, 1672448400, 1672452000, 1672455600, 1672459200, 
    1672462800, 1672466400, 1672470000, 1672473600, 1672477200, 1672480800, 
    1672484400, 1672488000, 1672491600, 1672495200, 1672498800, 1672502400, 
    1672506000, 1672509600, 1672513200, 1672516800, 1672520400, 1672524000, 
    1672527600 ;

 pressure_level = 1000, 925, 850, 700, 500, 200 ;

 latitude = 28, 27.75, 27.5, 27.25, 27, 26.75, 26.5, 26.25, 26, 25.75, 25.5, 
    25.25, 25, 24.75, 24.5, 24.25, 24, 23.75, 23.5, 23.25, 23, 22.75, 22.5, 
    22.25, 22, 21.75, 21.5, 21.25, 21, 20.75, 20.5, 20.25, 20, 19.75, 19.5, 
    19.25, 19 ;

 longitude = 109, 109.25, 109.5, 109.75, 110, 110.25, 110.5, 110.75, 111, 
    111.25, 111.5, 111.75, 112, 112.25, 112.5, 112.75, 113, 113.25, 113.5, 
    113.75, 114, 114.25, 114.5, 114.75, 115, 115.25, 115.5, 115.75, 116, 
    116.25, 116.5, 116.75, 117, 117.25, 117.5, 117.75, 118, 118.25, 118.5, 
    118.75, 119 ;

 expver = "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", 
    "0001", "0001", "0001", "0001" ;
}
