netcdf onedim {
dimensions:
	d1 = 1;
variables:
	char c;
	char c2(d1);
data:
  c = 'a';
  c2 = 'b';
}
