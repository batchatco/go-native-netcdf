netcdf test_multidim {
dimensions:
  time = 2 ;
  lat = 3 ;
  lon = 4 ;
  level = 5 ;

variables:
  // Coordinate variables (same name as dimension)
  double time(time) ;
    time:units = "hours since 2024-01-01" ;
    time:calendar = "standard" ;
  float lat(lat) ;
    lat:units = "degrees_north" ;
    lat:long_name = "latitude" ;
  float lon(lon) ;
    lon:units = "degrees_east" ;
    lon:long_name = "longitude" ;
  float level(level) ;
    level:units = "hPa" ;
    level:positive = "down" ;

  // 2D field
  float surface_temp(lat, lon) ;
    surface_temp:units = "K" ;
    surface_temp:long_name = "surface temperature" ;
    surface_temp:_FillValue = -999.0f ;

  // 3D field
  float air_temp(time, lat, lon) ;
    air_temp:units = "K" ;
    air_temp:long_name = "air temperature" ;

  // 4D field
  float wind_speed(time, level, lat, lon) ;
    wind_speed:units = "m/s" ;
    wind_speed:long_name = "wind speed" ;

  // 1D along different dimensions
  int time_step(time) ;
  short lat_index(lat) ;
  ubyte lon_flag(lon) ;

// global attributes:
  :Conventions = "CF-1.8" ;
  :title = "multi-dimensional test" ;
  :source = "synthetic data" ;

data:
  time = 0.0, 6.0 ;
  lat = -30.0, 0.0, 30.0 ;
  lon = -120.0, -60.0, 0.0, 60.0 ;
  level = 1000.0, 850.0, 700.0, 500.0, 300.0 ;

  surface_temp =
    300.1, 301.2, 302.3, 303.4,
    290.1, 291.2, 292.3, 293.4,
    280.1, 281.2, 282.3, 283.4 ;

  air_temp =
    300.0, 301.0, 302.0, 303.0,
    290.0, 291.0, 292.0, 293.0,
    280.0, 281.0, 282.0, 283.0,
    299.0, 300.0, 301.0, 302.0,
    289.0, 290.0, 291.0, 292.0,
    279.0, 280.0, 281.0, 282.0 ;

  wind_speed =
    10.1, 10.2, 10.3, 10.4,  10.5, 10.6, 10.7, 10.8,  10.9, 11.0, 11.1, 11.2,
    20.1, 20.2, 20.3, 20.4,  20.5, 20.6, 20.7, 20.8,  20.9, 21.0, 21.1, 21.2,
    30.1, 30.2, 30.3, 30.4,  30.5, 30.6, 30.7, 30.8,  30.9, 31.0, 31.1, 31.2,
    40.1, 40.2, 40.3, 40.4,  40.5, 40.6, 40.7, 40.8,  40.9, 41.0, 41.1, 41.2,
    50.1, 50.2, 50.3, 50.4,  50.5, 50.6, 50.7, 50.8,  50.9, 51.0, 51.1, 51.2,
    11.1, 11.2, 11.3, 11.4,  11.5, 11.6, 11.7, 11.8,  11.9, 12.0, 12.1, 12.2,
    21.1, 21.2, 21.3, 21.4,  21.5, 21.6, 21.7, 21.8,  21.9, 22.0, 22.1, 22.2,
    31.1, 31.2, 31.3, 31.4,  31.5, 31.6, 31.7, 31.8,  31.9, 32.0, 32.1, 32.2,
    41.1, 41.2, 41.3, 41.4,  41.5, 41.6, 41.7, 41.8,  41.9, 42.0, 42.1, 42.2,
    51.1, 51.2, 51.3, 51.4,  51.5, 51.6, 51.7, 51.8,  51.9, 52.0, 52.1, 52.2 ;

  time_step = 1, 2 ;
  lat_index = -1, 0, 1 ;
  lon_flag = 0, 1, 1, 0 ;
}
