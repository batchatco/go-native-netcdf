netcdf testvlen {
types:
  int(*) vint;
  compound Easy {
    int FirstEasy;
    int SecondEasy;
  };
  Easy(*) EasyVlen;
  compound Tricky_t {
    int TrickyInt;
    EasyVlen TrickVlen;
  };
dimensions:
  dim = 6;

variables:
  vint v(dim);
  Tricky_t v:Tricky = {1, {{2, 3}, {4, 5}, {6,7}}};

  vint v2(dim);
  vint v2:Vint = {}, {1}, {2,3}, {4,5,6}, {7,8,9,10}, {11,12,13,14,15};

  Tricky_t :Tricky = {1, {{2, 3}, {4, 5}, {6,7}}};
  vint :Vint = {}, {1}, {2,3}, {4,5,6}, {7,8,9,10}, {11,12,13,14,15};

data:
  v = {}, {1}, {2,3}, {4,5,6}, {7,8,9,10}, {11,12,13,14,15};
  v2 = {11,12,13,14,15}, {7,8,9,10}, {4,5,6}, {2,3}, {1}, {};
}
