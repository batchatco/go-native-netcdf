netcdf testempty {
types:
  opaque(5) opaque5;
  compound alltypes {
    byte b;
    short s;
    int i;
    float f;
    double d;
  };

dimensions:
        u = UNLIMITED ; // (0 currently)
variables:
        int a(u);
        opaque5 b(u);
        alltypes c(u);
        alltypes d(u,u);
        alltypes e(u,u,u);
        opaque5 f(u,u);
        opaque5 g(u,u,u);
data:
}
