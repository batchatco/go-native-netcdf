netcdf tst_mslp {
}
