netcdf testenum {
types:
  byte enum color {
    RED = 0,
    YELLOW = 1,
    GREEN = 2,
    CYAN = 3,
    BLUE = 4,
    MAGENTA = 5
  };
  ushort enum color2 {
    BLACK = 0,
    WHITE = 1
  };
  int64 enum junk {
    FIRST = 1L,
    SECOND = 2,
    THIRD = 3,
    FOURTH = 4,
    FIFTH = 5,
    SIXTH = 6
  };
  int enum junk2 {
    SEVENTH = 7,
    EIGHTH = 8
  };

dimensions:
  dim = 6;

variables:
  color nodim;
  color c(dim);
  junk j(dim);
  color2 c2;
  junk2 j2;

data:
  nodim = GREEN;

  c = RED, YELLOW, GREEN, CYAN, BLUE, MAGENTA;

  c2 = BLACK;

  j = FIRST, SECOND, THIRD, FOURTH, FIFTH, SIXTH;

  j2 = SEVENTH;
}
