netcdf testenum {
types:
  byte enum color {
    RED = 0,
    YELLOW = 1,
    GREEN = 2,
    CYAN = 3,
    BLUE = 4,
    MAGENTA = 5
  };
  int64 enum junk {
    FIRST = 1,
    SECOND = 2,
    THIRD = 3,
    FOURTH = 4,
    FIFTH = 5,
    SIXTH = 6
  };

dimensions:
  dim = 6;

variables:
  color nodim;
  color c(dim);
  junk j(dim);

data:
  nodim = GREEN;

  c = RED, YELLOW, GREEN, CYAN, BLUE, MAGENTA;

  j = FIRST, SECOND, THIRD, FOURTH, FIFTH, SIXTH;
}
