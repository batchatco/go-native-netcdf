netcdf testmultidim {
  dimensions:
	d1 = 2 ;
	d2 = 2 ;
	d3 = 3 ;
	d4 = 4 ;
variables:
	ushort val(d1, d2, d3, d4);
data:
  val =
    0, 1, 2, 3,
    4, 5, 6, 7,
    8, 9, 10, 11,
    12, 13, 14, 15,
    16, 17, 18, 19,
    20, 21, 22, 23,
    100, 101, 102, 103,
    104, 105, 106, 107,
    108, 109, 110, 111,
    112, 113, 114, 115,
    116, 117, 118, 119,
    120, 121, 122, 123;
}
