netcdf testnull {
}
