netcdf testempty {
dimensions:
  u = UNLIMITED ; // (0 currently)
variables:
  int a(u);
}
