netcdf testgroups {
dimensions:
  d1 = 1;
variables:
  int datamember(d1);
data:
  datamember = 2;
  group:  a {
    dimensions:
      d1 = 2;
    variables:
      int datamember(d1);
    data:
      datamember = 3, 4;

    group: b {
      dimensions:
        d1 = 3;
      variables:
        int datamember(d1);
      data:
        datamember = 5, 6, 7;
    }
  }
}
