netcdf testcompounds {
types:
  compound alltypes {
    byte b;
    short s;
    int i;
    float f;
    double d;
  };
  compound includes {
    alltypes a;
    string s;
  };
  compound sametypes {
    int a;
    int b;
    int c;
  };

dimensions:
  dim = UNLIMITED;

variables:
  includes v(dim);
  sametypes same(dim);

data:
  v = {{'0', 1, 2, 3.0, 4.0}, "a"}, {{'1', 2, 3, 4.0, 5.0}, "b"};

  same = {0,1,2},{3,4,5};
}
