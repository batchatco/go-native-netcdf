netcdf testslicer {
dimensions:
  lat = 4;
  lon = 5;
variables:
  byte tid(lat, lon);
data:
  tid = 0, 1, 2, 3, 4,
  5, 6, 6, 8, 9,
  10, 11, 12, 13, 14,
  15, 16, 17, 18, 19;
}
