netcdf testarray {
types:
	compound comp {
		int iArray(3);
		float fArray(2, 3);
	};
dimensions:
	dim = 2;
variables:
	comp c(dim);
data:
	c =
			{{1, 2, 3},
				{4, 5, 6, 7, 8, 9}},
			{{10, 11, 12},
				{13, 14, 15, 16, 17, 18}};
}
