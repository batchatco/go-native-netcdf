netcdf testunlimited {
dimensions:
	d1 = UNLIMITED;
variables:
	byte i8x1(d1);
data:
  i8x1 = 12, 56;
}
