netcdf filters {
dimensions:
  dim = 10;
variables:
  int nums(dim);
data:
  nums = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9;
}

