netcdf testvlen {
types:
  int(*) vint;

dimensions:
  dim = 5;

variables:
  vint v(dim);

data:
  v =  { 1 }, {2,3}, { 4,5,6}, {7,8,9,10},   {11,12,13,14,15};
}